
module bits ( clk, rst, pushin, datain, reqin, reqlen, pushout, lenout, 
        dataout );
  input [31:0] datain;
  input [3:0] reqlen;
  output [3:0] lenout;
  output [14:0] dataout;
  input clk, rst, pushin, reqin;
  output pushout;
  wire   pushin0, reqin0, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55,
         N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97,
         N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N310,
         N312, N313, N314, N317, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N436,
         N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448,
         N449, N450, N451, N452, N453, N456, N457, N458, N463, N465, N466,
         N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477,
         N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510,
         N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521,
         N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532,
         N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543,
         N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554,
         N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565,
         N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576,
         N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587,
         N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598,
         N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609,
         N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620,
         N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631,
         N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697,
         N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752,
         N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763,
         N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034,
         N1035, N1036, N1037, N1038, N1039, N1040, N1041, N2066, N2067, N2068,
         N2069, N2070, N2072, N2073, N2074, N2075, N2076, N2077, N2078, N2079,
         N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089,
         N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099,
         N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109,
         N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119,
         N2120, N2121, N2122, N2123, N2124, N2125, N2126, N2127, N2128, N2129,
         N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138, N2139,
         N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149,
         N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158, N2159,
         N2160, N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168, N2169,
         N2170, N2171, N2172, N2173, N2174, N2175, N2176, N2177, N2178, N2179,
         N2180, N2181, N2182, N2183, N2184, N2185, N2186, N2187, N2188, N2189,
         N2190, N2191, N2192, N2193, N2194, N2195, N2196, N2197, N2198, N2199,
         N2200, N2201, N2202, N2203, N2204, N2205, N2206, N2207, N2208, N2209,
         N2210, N2211, N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219,
         N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229,
         N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239,
         N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249,
         N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259,
         N2260, N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269,
         N2270, N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279,
         N2280, N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289,
         N2290, N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299,
         N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309,
         N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319,
         N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329,
         N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339,
         N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349,
         N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359,
         N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369,
         N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379,
         N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389,
         N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399,
         N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409,
         N2410, N2411, N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419,
         N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429,
         N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2438, N2439,
         N2440, N2441, N2442, N2443, N2444, N2445, N2446, N2447, N2448, N2449,
         N2450, N2451, N2452, N2453, N2454, N2455, N2456, N2457, N2458, N2459,
         N2460, N2461, N2462, N2463, N2464, N2465, N2466, N2467, N2468, N2469,
         N2470, N2471, N2472, N2473, N2474, N2475, N2476, N2477, N2478, N2479,
         N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489,
         N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499,
         N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509,
         N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519,
         N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529,
         N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539,
         N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, N2549,
         N2550, N2551, N2552, N2553, N2554, N2555, N2556, N2557, N2558, N2559,
         N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569,
         N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2579,
         N2580, N2581, N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589,
         N2590, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599,
         N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609,
         N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619,
         N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629,
         N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639,
         N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649,
         N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659,
         N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669,
         N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679,
         N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687, N2688, N2689,
         N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697, N2698, N2699,
         N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707, N2708, N2709,
         N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719,
         N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727, N2728, N2729,
         N2730, N2731, N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739,
         N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2749,
         N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757, N2758, N2759,
         N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769,
         N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779,
         N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789,
         N2790, N2791, N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799,
         N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809,
         N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819,
         N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829,
         N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839,
         N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849,
         N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859,
         N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869,
         N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879,
         N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889,
         N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899,
         N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909,
         N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919,
         N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929,
         N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939,
         N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949,
         N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959,
         N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969,
         N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979,
         N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989,
         N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999,
         N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009,
         N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019,
         N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029,
         N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039,
         N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049,
         N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059,
         N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069,
         N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079,
         N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089,
         N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099,
         N3105, N3106, N3107, N3108, N3109, N5158, N5159, N5160, N5161, N5162,
         N5163, N5164, N5165, N5166, N5167, N5168, N5169, N5170, N5171, N5172,
         N5173, N5174, N5175, N5176, N5177, N5178, N5179, N5180, N5181, N5182,
         N5183, N5184, N5185, N5186, N5187, N5188, N5189, N5190, N5191, N5192,
         N5193, N5194, N5195, N5196, N5197, N5198, N5199, N5200, N5201, N5202,
         N5203, N5204, N5205, N5206, N5207, N5208, N5209, N5210, N5211, N5212,
         N5213, N5214, N5215, N5216, N5217, N5218, N5219, N5220, N5221, N5222,
         N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5231, N5232,
         N5233, N5234, N5235, N5236, N5237, N5238, N5239, N5240, N5241, N5242,
         N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5251, N5252,
         N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262,
         N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271, N5272,
         N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281, N5282,
         N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291, N5292,
         N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5301, N5302,
         N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312,
         N5313, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321, N5322,
         N5323, N5324, N5325, N5326, N5327, N5328, N5329, N5330, N5331, N5332,
         N5333, N5334, N5335, N5336, N5337, N5338, N5339, N5340, N5341, N5342,
         N5343, N5344, N5345, N5346, N5347, N5348, N5349, N5350, N5351, N5352,
         N5353, N5354, N5355, N5356, N5357, N5358, N5359, N5360, N5361, N5362,
         N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5372,
         N5373, N5374, N5375, N5376, N5377, N5378, N5379, N5380, N5381, N5382,
         N5383, N5384, N5385, N5386, N5387, N5388, N5389, N5390, N5391, N5392,
         N5393, N5394, N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402,
         N5403, N5404, N5405, N5406, N5407, N5408, N5409, N5410, N5411, N5412,
         N5413, N5414, N5415, N5416, N5417, N5418, N5419, N5420, N5421, N5422,
         N5423, N5424, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5432,
         N5433, N5434, N5435, N5436, N5437, N5438, N5439, N5440, N5441, N5442,
         N5443, N5444, N5445, N5446, N5447, N5448, N5449, N5450, N5451, N5452,
         N5453, N5454, N5455, N5456, N5457, N5458, N5459, N5460, N5461, N5462,
         N5463, N5464, N5465, N5466, N5467, N5468, N5469, N5470, N5471, N5472,
         N5473, N5474, N5475, N5476, N5477, N5478, N5479, N5480, N5481, N5482,
         N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5490, N5491, N5492,
         N5493, N5494, N5495, N5496, N5497, N5498, N5499, N5500, N5501, N5502,
         N5503, N5504, N5505, N5506, N5507, N5508, N5509, N5510, N5511, N5512,
         N5513, N5514, N5515, N5516, N5517, N5518, N5519, N5520, N5521, N5522,
         N5523, N5524, N5525, N5526, N5527, N5528, N5529, N5530, N5531, N5532,
         N5533, N5534, N5535, N5536, N5537, N5538, N5539, N5540, N5541, N5542,
         N5543, N5544, N5545, N5546, N5547, N5548, N5549, N5550, N5551, N5552,
         N5553, N5554, N5555, N5556, N5557, N5558, N5559, N5560, N5561, N5562,
         N5563, N5564, N5565, N5566, N5567, N5568, N5569, N5570, N5571, N5572,
         N5573, N5574, N5575, N5576, N5577, N5578, N5579, N5580, N5581, N5582,
         N5583, N5584, N5585, N5586, N5587, N5588, N5589, N5590, N5591, N5592,
         N5593, N5594, N5595, N5596, N5597, N5598, N5599, N5600, N5601, N5602,
         N5603, N5604, N5605, N5606, N5607, N5608, N5609, N5610, N5611, N5612,
         N5613, N5614, N5615, N5616, N5617, N5618, N5619, N5620, N5621, N5622,
         N5623, N5624, N5625, N5626, N5627, N5628, N5629, N5630, N5631, N5632,
         N5633, N5634, N5635, N5636, N5637, N5638, N5639, N5640, N5641, N5642,
         N5643, N5644, N5645, N5646, N5647, N5648, N5649, N5650, N5651, N5652,
         N5653, N5654, N5655, N5656, N5657, N5658, N5659, N5660, N5661, N5662,
         N5663, N5664, N5665, N5666, N5667, N5668, N5669, N5670, N5671, N5672,
         N5673, N5674, N5675, N5676, N5677, N5678, N5679, N5680, N5681, N5682,
         N5683, N5684, N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692,
         N5693, N5694, N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702,
         N5703, N5704, N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712,
         N5713, N5714, N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722,
         N5723, N5724, N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732,
         N5733, N5734, N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742,
         N5743, N5744, N5745, N5746, N5747, N5748, N5749, N5750, N5751, N5752,
         N5753, N5754, N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762,
         N5763, N5764, N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772,
         N5773, N5774, N5775, N5776, N5777, N5778, N5779, N5780, N5781, N5782,
         N5783, N5784, N5785, N5786, N5787, N5788, N5789, N5790, N5791, N5792,
         N5793, N5794, N5795, N5796, N5797, N5798, N5799, N5800, N5801, N5802,
         N5803, N5804, N5805, N5806, N5807, N5808, N5809, N5810, N5811, N5812,
         N5813, N5814, N5815, N5816, N5817, N5818, N5819, N5820, N5821, N5822,
         N5823, N5824, N5825, N5826, N5827, N5828, N5829, N5830, N5831, N5832,
         N5833, N5834, N5835, N5836, N5837, N5838, N5839, N5840, N5841, N5842,
         N5843, N5844, N5845, N5846, N5847, N5848, N5849, N5850, N5851, N5852,
         N5853, N5854, N5855, N5856, N5857, N5858, N5859, N5860, N5861, N5862,
         N5863, N5864, N5865, N5866, N5867, N5868, N5869, N5870, N5871, N5872,
         N5873, N5874, N5875, N5876, N5877, N5878, N5879, N5880, N5881, N5882,
         N5883, N5884, N5885, N5886, N5887, N5888, N5889, N5890, N5891, N5892,
         N5893, N5894, N5895, N5896, N5897, N5898, N5899, N5900, N5901, N5902,
         N5903, N5904, N5905, N5906, N5907, N5908, N5909, N5910, N5911, N5912,
         N5913, N5914, N5915, N5916, N5917, N5918, N5919, N5920, N5921, N5922,
         N5923, N5924, N5925, N5926, N5927, N5928, N5929, N5930, N5931, N5932,
         N5933, N5934, N5935, N5936, N5937, N5938, N5939, N5940, N5941, N5942,
         N5943, N5944, N5945, N5946, N5947, N5948, N5949, N5950, N5951, N5952,
         N5953, N5954, N5955, N5956, N5957, N5958, N5959, N5960, N5961, N5962,
         N5963, N5964, N5965, N5966, N5967, N5968, N5969, N5970, N5971, N5972,
         N5973, N5974, N5975, N5976, N5977, N5978, N5979, N5980, N5981, N5982,
         N5983, N5984, N5985, N5986, N5987, N5988, N5989, N5990, N5991, N5992,
         N5993, N5994, N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002,
         N6003, N6004, N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012,
         N6013, N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022,
         N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032,
         N6033, N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6042,
         N6043, N6044, N6045, N6046, N6047, N6048, N6049, N6050, N6051, N6052,
         N6053, N6054, N6055, N6056, N6057, N6058, N6059, N6060, N6061, N6062,
         N6063, N6064, N6065, N6066, N6067, N6068, N6069, N6070, N6071, N6072,
         N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6081, N6082,
         N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6092,
         N6093, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102,
         N6103, N6104, N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112,
         N6113, N6114, N6115, N6116, N6117, N6118, N6119, N6120, N6121, N6122,
         N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132,
         N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6141, N6142,
         N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6150, N6151, N6152,
         N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162,
         N6163, N6164, N6165, N6166, N6167, N6168, N6169, N6170, N6171, N6172,
         N6173, N6174, N6175, N6176, N6177, N6178, N6179, N6180, N6181, N6222,
         N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231, N7256,
         N7257, N7258, N7259, N7260, N7261, N7262, N7263, N7264, N7265, N7266,
         N7267, N7268, N7269, N7270, N7271, N7272, N7273, N7274, N7275, N7276,
         N7277, N7278, N7279, N7280, N7281, N7282, N7283, N7284, N7285, N7286,
         N7287, N7288, N7289, N7290, N7291, N7292, N7293, N7294, N7295, N7296,
         N7297, N7298, N7299, N7300, N7301, N7302, N7303, N7304, N7305, N7306,
         N7307, N7308, N7309, N7310, N7311, N7312, N7313, N7314, N7315, N7316,
         N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7325, N7326,
         N7327, N7328, N7329, N7330, N7331, N7332, N7333, N7334, N7335, N7336,
         N7337, N7338, N7339, N7340, N7341, N7342, N7343, N7344, N7345, N7346,
         N7347, N7348, N7349, N7350, N7351, N7352, N7353, N7354, N7355, N7356,
         N7357, N7358, N7359, N7360, N7361, N7362, N7363, N7364, N7365, N7366,
         N7367, N7368, N7369, N7370, N7371, N7372, N7373, N7374, N7375, N7376,
         N7377, N7378, N7379, N7380, N7381, N7382, N7383, N7384, N7385, N7386,
         N7387, N7388, N7389, N7390, N7391, N7392, N7393, N7394, N7395, N7396,
         N7397, N7398, N7399, N7400, N7401, N7402, N7403, N7404, N7405, N7406,
         N7407, N7408, N7409, N7410, N7411, N7412, N7413, N7414, N7415, N7416,
         N7417, N7418, N7419, N7420, N7421, N7422, N7423, N7424, N7425, N7426,
         N7427, N7428, N7429, N7430, N7431, N7432, N7433, N7434, N7435, N7436,
         N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446,
         N7447, N7448, N7449, N7450, N7451, N7452, N7453, N7454, N7455, N7456,
         N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7465, N7466,
         N7467, N7468, N7469, N7470, N7471, N7472, N7473, N7474, N7475, N7476,
         N7477, N7478, N7479, N7480, N7481, N7482, N7483, N7484, N7485, N7486,
         N7487, N7488, N7489, N7490, N7491, N7492, N7493, N7494, N7495, N7496,
         N7497, N7498, N7499, N7500, N7501, N7502, N7503, N7504, N7505, N7506,
         N7507, N7508, N7509, N7510, N7511, N7512, N7513, N7514, N7515, N7516,
         N7517, N7518, N7519, N7520, N7521, N7522, N7523, N7524, N7525, N7526,
         N7527, N7528, N7529, N7530, N7531, N7532, N7533, N7534, N7535, N7536,
         N7537, N7538, N7539, N7540, N7541, N7542, N7543, N7544, N7545, N7546,
         N7547, N7548, N7549, N7550, N7551, N7552, N7553, N7554, N7555, N7556,
         N7557, N7558, N7559, N7560, N7561, N7562, N7563, N7564, N7565, N7566,
         N7567, N7568, N7569, N7570, N7571, N7572, N7573, N7574, N7575, N7576,
         N7577, N7578, N7579, N7580, N7581, N7582, N7583, N7584, N7585, N7586,
         N7587, N7588, N7589, N7590, N7591, N7592, N7593, N7594, N7595, N7596,
         N7597, N7598, N7599, N7600, N7601, N7602, N7603, N7604, N7605, N7606,
         N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, N7615, N7616,
         N7617, N7618, N7619, N7620, N7621, N7622, N7623, N7624, N7625, N7626,
         N7627, N7628, N7629, N7630, N7631, N7632, N7633, N7634, N7635, N7636,
         N7637, N7638, N7639, N7640, N7641, N7642, N7643, N7644, N7645, N7646,
         N7647, N7648, N7649, N7650, N7651, N7652, N7653, N7654, N7655, N7656,
         N7657, N7658, N7659, N7660, N7661, N7662, N7663, N7664, N7665, N7666,
         N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676,
         N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686,
         N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696,
         N7697, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7708, N7709, N7710, N7711, N7712, N7713, N7714, N7715, N7716,
         N7717, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7725, N7726,
         N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7735, N7736,
         N7737, N7738, N7739, N7740, N7741, N7742, N7743, N7744, N7745, N7746,
         N7747, N7748, N7749, N7750, N7751, N7752, N7753, N7754, N7755, N7756,
         N7757, N7758, N7759, N7760, N7761, N7762, N7763, N7764, N7765, N7766,
         N7767, N7768, N7769, N7770, N7771, N7772, N7773, N7774, N7775, N7776,
         N7777, N7778, N7779, N7780, N7781, N7782, N7783, N7784, N7785, N7786,
         N7787, N7788, N7789, N7790, N7791, N7792, N7793, N7794, N7795, N7796,
         N7797, N7798, N7799, N7800, N7801, N7802, N7803, N7804, N7805, N7806,
         N7807, N7808, N7809, N7810, N7811, N7812, N7813, N7814, N7815, N7816,
         N7817, N7818, N7819, N7820, N7821, N7822, N7823, N7824, N7825, N7826,
         N7827, N7828, N7829, N7830, N7831, N7832, N7833, N7834, N7835, N7836,
         N7837, N7838, N7839, N7840, N7841, N7842, N7843, N7844, N7845, N7846,
         N7847, N7848, N7849, N7850, N7851, N7852, N7853, N7854, N7855, N7856,
         N7857, N7858, N7859, N7860, N7861, N7862, N7863, N7864, N7865, N7866,
         N7867, N7868, N7869, N7870, N7871, N7872, N7873, N7874, N7875, N7876,
         N7877, N7878, N7879, N7880, N7881, N7882, N7883, N7884, N7885, N7886,
         N7887, N7888, N7889, N7890, N7891, N7892, N7893, N7894, N7895, N7896,
         N7897, N7898, N7899, N7900, N7901, N7902, N7903, N7904, N7905, N7906,
         N7907, N7908, N7909, N7910, N7911, N7912, N7913, N7914, N7915, N7916,
         N7917, N7918, N7919, N7920, N7921, N7922, N7923, N7924, N7925, N7926,
         N7927, N7928, N7929, N7930, N7931, N7932, N7933, N7934, N7935, N7936,
         N7937, N7938, N7939, N7940, N7941, N7942, N7943, N7944, N7945, N7946,
         N7947, N7948, N7949, N7950, N7951, N7952, N7953, N7954, N7955, N7956,
         N7957, N7958, N7959, N7960, N7961, N7962, N7963, N7964, N7965, N7966,
         N7967, N7968, N7969, N7970, N7971, N7972, N7973, N7974, N7975, N7976,
         N7977, N7978, N7979, N7980, N7981, N7982, N7983, N7984, N7985, N7986,
         N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996,
         N7997, N7998, N7999, N8000, N8001, N8002, N8003, N8004, N8005, N8006,
         N8007, N8008, N8009, N8010, N8011, N8012, N8013, N8014, N8015, N8016,
         N8017, N8018, N8019, N8020, N8021, N8022, N8023, N8024, N8025, N8026,
         N8027, N8028, N8029, N8030, N8031, N8032, N8033, N8034, N8035, N8036,
         N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8046,
         N8047, N8048, N8049, N8050, N8051, N8052, N8053, N8054, N8055, N8056,
         N8057, N8058, N8059, N8060, N8061, N8062, N8063, N8064, N8065, N8066,
         N8067, N8068, N8069, N8070, N8071, N8072, N8073, N8074, N8075, N8076,
         N8077, N8078, N8079, N8080, N8081, N8082, N8083, N8084, N8085, N8086,
         N8087, N8088, N8089, N8090, N8091, N8092, N8093, N8094, N8095, N8096,
         N8097, N8098, N8099, N8100, N8101, N8102, N8103, N8104, N8105, N8106,
         N8107, N8108, N8109, N8110, N8111, N8112, N8113, N8114, N8115, N8116,
         N8117, N8118, N8119, N8120, N8121, N8122, N8123, N8124, N8125, N8126,
         N8127, N8128, N8129, N8130, N8131, N8132, N8133, N8134, N8135, N8136,
         N8137, N8138, N8139, N8140, N8141, N8142, N8143, N8144, N8145, N8146,
         N8147, N8148, N8149, N8150, N8151, N8152, N8153, N8154, N8155, N8156,
         N8157, N8158, N8159, N8160, N8161, N8162, N8163, N8164, N8165, N8166,
         N8167, N8168, N8169, N8170, N8171, N8172, N8173, N8174, N8175, N8176,
         N8177, N8178, N8179, N8180, N8181, N8182, N8183, N8184, N8185, N8186,
         N8187, N8188, N8189, N8190, N8191, N8192, N8193, N8194, N8195, N8196,
         N8197, N8198, N8199, N8200, N8201, N8202, N8203, N8204, N8205, N8206,
         N8207, N8208, N8209, N8210, N8211, N8212, N8213, N8214, N8215, N8216,
         N8217, N8218, N8219, N8220, N8221, N8222, N8223, N8224, N8225, N8226,
         N8227, N8228, N8229, N8230, N8231, N8232, N8233, N8234, N8235, N8236,
         N8237, N8238, N8239, N8240, N8241, N8242, N8243, N8244, N8245, N8246,
         N8247, N8248, N8249, N8250, N8251, N8252, N8253, N8254, N8255, N8256,
         N8257, N8258, N8259, N8260, N8261, N8262, N8263, N8264, N8265, N8266,
         N8267, N8268, N8269, N8270, N8271, N8272, N8273, N8274, N8275, N8276,
         N8277, N8278, N8279, N8280, N8281, N8282, N8283, N8284, N8285, N8286,
         N8287, N8288, N8289, N8290, N8291, N8292, N8293, N8294, N8295, N8296,
         N8297, N8298, N8299, N8300, N8301, N8302, N8303, N8304, N8305, N8306,
         N8307, N8308, N8309, N8310, N8311, N8312, N8313, N8314, N8315, N8316,
         N8317, N8318, N8319, N8320, N8321, N8322, N8323, N8324, N8325, N8326,
         N8327, N8328, N8329, N8330, N8331, N8332, N8333, N8334, N8335, N8336,
         N8337, N8338, N8339, N8340, N8341, N8342, N8343, N8344, N8345, N8346,
         N8347, N8348, N8349, N8350, N8351, N8352, N8353, N8354, N8355, N8356,
         N8357, N8358, N8359, N8360, N8361, N8362, N8363, N8364, N8365, N8366,
         N8367, N8368, N8369, N8370, N8371, N8372, N8373, N8374, N8375, N8376,
         N8377, N8378, N8379, N8380, N8381, N8382, N8383, N8384, N8385, N8386,
         N8387, N8388, N8389, N8390, N8391, N8392, N8393, N8394, N8395, N8396,
         N8397, N8398, N8399, N8400, N8401, N8402, N8403, N8404, N8405, N8406,
         N8407, N8408, N8409, N8410, N8411, N8412, N8413, N8414, N8415, N8416,
         N8417, N8418, N8419, N8420, N8421, N8422, N8423, N8424, N8425, N8426,
         N8427, N8428, N8429, N8430, N8431, N8432, N8433, N8434, N8435, N8436,
         N8437, N8438, N8439, N8440, N8441, N8442, N8443, N8444, N8445, N8446,
         N8447, N8448, N8449, N8450, N8451, N8452, N8453, N8454, N8455, N8456,
         N8457, N8458, N8459, N8460, N8461, N8462, N8463, N8464, N8465, N8466,
         N8467, N8468, N8469, N8470, N8471, N8472, N8473, N8474, N8475, N8476,
         N8477, N8478, N8479, N8480, N8481, N8482, N8483, N8484, N8485, N8486,
         N8487, N8488, N8489, N8490, N8491, N8492, N8493, N8494, N8495, N8496,
         N8497, N8498, N8499, N8500, N8501, N8502, N8503, N8504, N8505, N8506,
         N8507, N8508, N8509, N8510, N8511, N8512, N8513, N8514, N8515, N8516,
         N8517, N8518, N8519, N8520, N8521, N8522, N8523, N8524, N8525, N8526,
         N8527, N8528, N8529, N8530, N8531, N8532, N8533, N8534, N8535, N8536,
         N8537, N8538, N8539, N8540, N8541, N8542, N8543, N8544, N8545, N8546,
         N8547, N8548, N8549, N8550, N8551, N8552, N8553, N8554, N8555, N8556,
         N8557, N8558, N8559, N8560, N8561, N8562, N8563, N8564, N8565, N8566,
         N8567, N8568, N8569, N8570, N8571, N8572, N8573, N8574, N8575, N8576,
         N8577, N8578, N8579, N8580, N8581, N8582, N8583, N8584, N8585, N8586,
         N8587, N8588, N8589, N8590, N8591, N8592, N8593, N8594, N8595, N8596,
         N8597, N8598, N8599, N8600, N8601, N8602, N8603, N8604, N8605, N8606,
         N8607, N8608, N8609, N8610, N8611, N8612, N8613, N8614, N8615, N8616,
         N8617, N8618, N8619, N8620, N8621, N8622, N8623, N8624, N8625, N8626,
         N8627, N8628, N8629, N8630, N8631, N8632, N8633, N8634, N8635, N8636,
         N8637, N8638, N8639, N8640, N8641, N8642, N8643, N8644, N8645, N8646,
         N8647, N8648, N8649, N8650, N8651, N8652, N8653, N8654, N8655, N8656,
         N8657, N8658, N8659, N8660, N8661, N8662, N8663, N8664, N8665, N8666,
         N8667, N8668, N8669, N8670, N8671, N8672, N8673, N8674, N8675, N8676,
         N8677, N8678, N8679, N8680, N8681, N8682, N8683, N8684, N8685, N8686,
         N8687, N8688, N8689, N8690, N8691, N8692, N8693, N8694, N8695, N8696,
         N8697, N8698, N8699, N8700, N8701, N8702, N8703, N8704, N8705, N8706,
         N8707, N8708, N8709, N8710, N8711, N8712, N8713, N8714, N8715, N8716,
         N8717, N8718, N8719, N8720, N8721, N8722, N8723, N8724, N8725, N8726,
         N8727, N8728, N8729, N8730, N8731, N8732, N8733, N8734, N8735, N8736,
         N8737, N8738, N8739, N8740, N8741, N8742, N8743, N8744, N8745, N8746,
         N8747, N8748, N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756,
         N8757, N8758, N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766,
         N8767, N8768, N8769, N8770, N8771, N8772, N8773, N8774, N8775, N8776,
         N8777, N8778, N8779, N8780, N8781, N8782, N8783, N8784, N8785, N8786,
         N8787, N8788, N8789, N8790, N8791, N8792, N8793, N8794, N8795, N8796,
         N8797, N8798, N8799, N8800, N8801, N8802, N8803, N8804, N8805, N8806,
         N8807, N8808, N8809, N8810, N8811, N8812, N8813, N8814, N8815, N8816,
         N8817, N8818, N8819, N8820, N8821, N8822, N8823, N8824, N8825, N8826,
         N8827, N8828, N8829, N8830, N8831, N8832, N8833, N8834, N8835, N8836,
         N8837, N8838, N8839, N8840, N8841, N8842, N8843, N8844, N8845, N8846,
         N8847, N8848, N8849, N8850, N8851, N8852, N8853, N8854, N8855, N8856,
         N8857, N8858, N8859, N8860, N8861, N8862, N8863, N8864, N8865, N8866,
         N8867, N8868, N8869, N8870, N8871, N8872, N8873, N8874, N8875, N8876,
         N8877, N8878, N8879, N8880, N8881, N8882, N8883, N8884, N8885, N8886,
         N8887, N8888, N8889, N8890, N8891, N8892, N8893, N8894, N8895, N8896,
         N8897, N8898, N8899, N8900, N8901, N8902, N8903, N8904, N8905, N8906,
         N8907, N8908, N8909, N8910, N8911, N8912, N8913, N8914, N8915, N8916,
         N8917, N8918, N8919, N8920, N8921, N8922, N8923, N8924, N8925, N8926,
         N8927, N8928, N8929, N8930, N8931, N8932, N8933, N8934, N8935, N8936,
         N8937, N8938, N8939, N8940, N8941, N8942, N8943, N8944, N8945, N8946,
         N8947, N8948, N8949, N8950, N8951, N8952, N8953, N8954, N8955, N8956,
         N8957, N8958, N8959, N8960, N8961, N8962, N8963, N8964, N8965, N8966,
         N8967, N8968, N8969, N8970, N8971, N8972, N8973, N8974, N8975, N8976,
         N8977, N8978, N8979, N8980, N8981, N8982, N8983, N8984, N8985, N8986,
         N8987, N8988, N8989, N8990, N8991, N8992, N8993, N8994, N8995, N8996,
         N8997, N8998, N8999, N9000, N9001, N9002, N9003, N9004, N9005, N9006,
         N9007, N9008, N9009, N9010, N9011, N9012, N9013, N9014, N9015, N9016,
         N9017, N9018, N9019, N9020, N9021, N9022, N9023, N9024, N9025, N9026,
         N9027, N9028, N9029, N9030, N9031, N9032, N9033, N9034, N9035, N9036,
         N9037, N9038, N9039, N9040, N9041, N9042, N9043, N9044, N9045, N9046,
         N9047, N9048, N9049, N9050, N9051, N9052, N9053, N9054, N9055, N9056,
         N9057, N9058, N9059, N9060, N9061, N9062, N9063, N9064, N9065, N9066,
         N9067, N9068, N9069, N9070, N9071, N9072, N9073, N9074, N9075, N9076,
         N9077, N9078, N9079, N9080, N9081, N9082, N9083, N9084, N9085, N9086,
         N9087, N9088, N9089, N9090, N9091, N9092, N9093, N9094, N9095, N9096,
         N9097, N9098, N9099, N9100, N9101, N9102, N9103, N9104, N9105, N9106,
         N9107, N9108, N9109, N9110, N9111, N9112, N9113, N9114, N9115, N9116,
         N9117, N9118, N9119, N9120, N9121, N9122, N9123, N9124, N9125, N9126,
         N9127, N9128, N9129, N9130, N9131, N9132, N9133, N9134, N9135, N9136,
         N9137, N9138, N9139, N9140, N9141, N9142, N9143, N9144, N9145, N9146,
         N9147, N9148, N9149, N9150, N9151, N9152, N9153, N9154, N9155, N9156,
         N9157, N9158, N9159, N9160, N9161, N9162, N9163, N9164, N9165, N9166,
         N9167, N9168, N9169, N9170, N9171, N9172, N9173, N9174, N9175, N9176,
         N9177, N9178, N9179, N9180, N9181, N9182, N9183, N9184, N9185, N9186,
         N9187, N9188, N9189, N9190, N9191, N9192, N9193, N9194, N9195, N9196,
         N9197, N9198, N9199, N9200, N9201, N9202, N9203, N9204, N9205, N9206,
         N9207, N9208, N9209, N9210, N9211, N9212, N9213, N9214, N9215, N9216,
         N9217, N9218, N9219, N9220, N9221, N9222, N9223, N9224, N9225, N9226,
         N9227, N9228, N9229, N9230, N9231, N9232, N9233, N9234, N9235, N9236,
         N9237, N9238, N9239, N9240, N9241, N9242, N9243, N9244, N9245, N9246,
         N9247, N9248, N9249, N9250, N9251, N9252, N9253, N9254, N9255, N9256,
         N9257, N9258, N9259, N9260, N9261, N9262, N9263, N9264, N9265, N9266,
         N9267, N9268, N9269, N9270, N9271, N9272, N9273, N9274, N9275, N9276,
         N9277, N9278, N9279, N9280, N9281, N9282, N9283, N9284, N9285, N9286,
         N9287, N9288, N9289, N9290, N9291, N9292, N9293, N9294, N9295, N9296,
         N9297, N9298, N9299, N9300, N9301, N9302, N9303, N9324, N9325, N9326,
         N9327, N9328, N9329, N9330, N9331, N9332, N9333, N9334, N9335, N9336,
         N9337, N9338, N9339, N9340, N9341, N9342, N9343, N9344, N9345, N9346,
         N9347, N9348, N9349, N9350, N9351, N9352, N9353, N9354, N9355, N9356,
         N9357, N9358, N9359, N9360, N9361, N9362, N9363, N9364, N9365, N9366,
         N9367, N9368, N9369, N9370, N9371, N9372, N9373, N9374, N9375, N9376,
         N9377, N9378, N9379, N9380, N9381, N9382, N9383, N9384, N9385, N9386,
         N9387, N9388, N9389, N9390, N9391, N9392, N9393, N9394, N9395, N9396,
         N9397, N9398, N9399, N9400, N9401, N9402, N9403, N9404, N9405, N9406,
         N9407, N9408, N9409, N9410, N9411, N9412, N9413, N9414, N9415, N9416,
         N9417, N9418, N9419, N9420, N9421, N9422, N9423, N9424, N9425, N9426,
         N9427, N9428, N9429, N9430, N9431, N9432, N9433, N9434, N9435, N9436,
         N9437, N9438, N9439, N9440, N9441, N9442, N9443, N9444, N9445, N9446,
         N9447, N9448, N9449, N9450, N9451, N9452, N9453, N9454, N9455, N9456,
         N9457, N9458, N9459, N9460, N9461, N9462, N9463, N9464, N9465, N9466,
         N9467, N9468, N9469, N9470, N9471, N9472, N9473, N9474, N9475, N9476,
         N9477, N9478, N9479, N9480, N9481, N9482, N9483, N9484, N9485, N9486,
         N9487, N9488, N9489, N9490, N9491, N9492, N9493, N9494, N9495, N9496,
         N9497, N9498, N9499, N9500, N9501, N9502, N9503, N9504, N9505, N9506,
         N9507, N9508, N9509, N9510, N9511, N9512, N9513, N9514, N9515, N9516,
         N9517, N9518, N9519, N9520, N9521, N9522, N9523, N9524, N9525, N9526,
         N9527, N9528, N9529, N9530, N9531, N9532, N9533, N9534, N9535, N9536,
         N9537, N9538, N9539, N9540, N9541, N9542, N9543, N9544, N9545, N9546,
         N9547, N9548, N9549, N9550, N9551, N9552, N9553, N9554, N9555, N9556,
         N9557, N9558, N9559, N9560, N9561, N9562, N9563, N9564, N9565, N9566,
         N9567, N9568, N9569, N9570, N9571, N9572, N9573, N9574, N9575, N9576,
         N9577, N9578, N9579, N9580, N9581, N9582, N9583, N9584, N9585, N9586,
         N9587, N9588, N9589, N9590, N9591, N9592, N9593, N9594, N9595, N9596,
         N9597, N9598, N9599, N9600, N9601, N9602, N9603, N9604, N9605, N9606,
         N9607, N9608, N9609, N9610, N9611, N9612, N9613, N9614, N9615, N9616,
         N9617, N9618, N9619, N9620, N9621, N9622, N9623, N9624, N9625, N9626,
         N9627, N9628, N9629, N9630, N9631, N9632, N9633, N9634, N9635, N9636,
         N9637, N9638, N9639, N9640, N9641, N9642, N9643, N9644, N9645, N9646,
         N9647, N9648, N9649, N9650, N9651, N9652, N9653, N9654, N9655, N9656,
         N9657, N9658, N9659, N9660, N9661, N9662, N9663, N9664, N9665, N9666,
         N9667, N9668, N9669, N9670, N9671, N9672, N9673, N9674, N9675, N9676,
         N9677, N9678, N9679, N9680, N9681, N9682, N9683, N9684, N9685, N9686,
         N9687, N9688, N9689, N9690, N9691, N9692, N9693, N9694, N9695, N9696,
         N9697, N9698, N9699, N9700, N9701, N9702, N9703, N9704, N9705, N9706,
         N9707, N9708, N9709, N9710, N9711, N9712, N9713, N9714, N9715, N9716,
         N9717, N9718, N9719, N9720, N9721, N9722, N9723, N9724, N9725, N9726,
         N9727, N9728, N9729, N9730, N9731, N9732, N9733, N9734, N9735, N9736,
         N9737, N9738, N9739, N9740, N9741, N9742, N9743, N9744, N9745, N9746,
         N9747, N9748, N9749, N9750, N9751, N9752, N9753, N9754, N9755, N9756,
         N9757, N9758, N9759, N9760, N9761, N9762, N9763, N9764, N9765, N9766,
         N9767, N9768, N9769, N9770, N9771, N9772, N9773, N9774, N9775, N9776,
         N9777, N9778, N9779, N9780, N9781, N9782, N9783, N9784, N9785, N9786,
         N9787, N9788, N9789, N9790, N9791, N9792, N9793, N9794, N9795, N9796,
         N9797, N9798, N9799, N9800, N9801, N9802, N9803, N9804, N9805, N9806,
         N9807, N9808, N9809, N9810, N9811, N9812, N9813, N9814, N9815, N9816,
         N9817, N9818, N9819, N9820, N9821, N9822, N9823, N9824, N9825, N9826,
         N9827, N9828, N9829, N9830, N9831, N9832, N9833, N9834, N9835, N9836,
         N9837, N9838, N9839, N9840, N9841, N9842, N9843, N9844, N9845, N9846,
         N9847, N9848, N9849, N9850, N9851, N9852, N9853, N9854, N9855, N9856,
         N9857, N9858, N9859, N9860, N9861, N9862, N9863, N9864, N9865, N9866,
         N9867, N9868, N9869, N9870, N9871, N9872, N9873, N9874, N9875, N9876,
         N9877, N9878, N9879, N9880, N9881, N9882, N9883, N9884, N9885, N9886,
         N9887, N9888, N9889, N9890, N9891, N9892, N9893, N9894, N9895, N9896,
         N9897, N9898, N9899, N9900, N9901, N9902, N9903, N9904, N9905, N9906,
         N9907, N9908, N9909, N9910, N9911, N9912, N9913, N9914, N9915, N9916,
         N9917, N9918, N9919, N9920, N9921, N9922, N9923, N9924, N9925, N9926,
         N9927, N9928, N9929, N9930, N9931, N9932, N9933, N9934, N9935, N9936,
         N9937, N9938, N9939, N9940, N9941, N9942, N9943, N9944, N9945, N9946,
         N9947, N9948, N9949, N9950, N9951, N9952, N9953, N9954, N9955, N9956,
         N9957, N9958, N9959, N9960, N9961, N9962, N9963, N9964, N9965, N9966,
         N9967, N9968, N9969, N9970, N9971, N9972, N9973, N9974, N9975, N9976,
         N9977, N9978, N9979, N9980, N9981, N9982, N9983, N9984, N9985, N9986,
         N9987, N9988, N9989, N9990, N9991, N9992, N9993, N9994, N9995, N9996,
         N9997, N9998, N9999, N10000, N10001, N10002, N10003, N10004, N10005,
         N10006, N10007, N10008, N10009, N10010, N10011, N10012, N10013,
         N10014, N10015, N10016, N10017, N10018, N10019, N10020, N10021,
         N10022, N10023, N10024, N10025, N10026, N10027, N10028, N10029,
         N10030, N10031, N10032, N10033, N10034, N10035, N10036, N10037,
         N10038, N10039, N10040, N10041, N10042, N10043, N10044, N10045,
         N10046, N10047, N10048, N10049, N10050, N10051, N10052, N10053,
         N10054, N10055, N10056, N10057, N10058, N10059, N10060, N10061,
         N10062, N10063, N10064, N10065, N10066, N10067, N10068, N10069,
         N10070, N10071, N10072, N10073, N10074, N10075, N10076, N10077,
         N10078, N10079, N10080, N10081, N10082, N10083, N10084, N10085,
         N10086, N10087, N10088, N10089, N10090, N10091, N10092, N10093,
         N10094, N10095, N10096, N10097, N10098, N10099, N10100, N10101,
         N10102, N10103, N10104, N10105, N10106, N10107, N10108, N10109,
         N10110, N10111, N10112, N10113, N10114, N10115, N10116, N10117,
         N10118, N10119, N10120, N10121, N10122, N10123, N10124, N10125,
         N10126, N10127, N10128, N10129, N10130, N10131, N10132, N10133,
         N10134, N10135, N10136, N10137, N10138, N10139, N10140, N10141,
         N10142, N10143, N10144, N10145, N10146, N10147, N10148, N10149,
         N10150, N10151, N10152, N10153, N10154, N10155, N10156, N10157,
         N10158, N10159, N10160, N10161, N10162, N10163, N10164, N10165,
         N10166, N10167, N10168, N10169, N10170, N10171, N10172, N10173,
         N10174, N10175, N10176, N10177, N10178, N10179, N10180, N10181,
         N10182, N10183, N10184, N10185, N10186, N10187, N10188, N10189,
         N10190, N10191, N10192, N10193, N10194, N10195, N10196, N10197,
         N10198, N10199, N10200, N10201, N10202, N10203, N10204, N10205,
         N10206, N10207, N10208, N10209, N10210, N10211, N10212, N10213,
         N10214, N10215, N10216, N10217, N10218, N10219, N10220, N10221,
         N10222, N10223, N10224, N10225, N10226, N10227, N10228, N10229,
         N10230, N10231, N10232, N10233, N10234, N10235, N10236, N10237,
         N10238, N10239, N10240, N10241, N10242, N10243, N10244, N10245,
         N10246, N10247, N10248, N10249, N10250, N10251, N10252, N10253,
         N10254, N10255, N10256, N10257, N10258, N10259, N10260, N10261,
         N10262, N10263, N10264, N10265, N10266, N10267, N10268, N10269,
         N10270, N10271, N10272, N10273, N10274, N10275, N10276, N10277,
         N10278, N10279, N10280, N10281, N10282, N10283, N10284, N10285,
         N10286, N10287, N10288, N10289, N10290, N10291, N10292, N10293,
         N10294, N10295, N10296, N10297, N10298, N10299, N10300, N10301,
         N10302, N10303, N10304, N10305, N10306, N10307, N10308, N10309,
         N10310, N10311, N10312, N10313, N10314, N10315, N10316, N10317,
         N10318, N10319, N10320, N10321, N10322, N10323, N10324, N10325,
         N10326, N10327, N10328, N10329, N10330, N10331, N10332, N10333,
         N10334, N10335, N10336, N10337, N10338, N10339, N10340, N10341,
         N10342, N10343, N10344, N10345, N10346, N10347, N10348, N10349,
         N10350, N10351, N10352, N10353, N10354, N10355, N10356, N10357,
         N10358, N10376, N10377, N10378, N10379, N10380, N10381, N10382,
         N10384, N10385, N10386, N10387, N10388, N10389, N10390, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n55,
         n56, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738;
  wire   [9:0] wr_ptr;
  wire   [3:0] lenin0;
  wire   [31:0] datain0;
  wire   [1023:0] mem_data1;
  wire   [10:0] \sub_84/carry ;
  wire   [10:0] \r349/carry ;
  wire   [9:1] \r347/carry ;

  COR2X1 U5218 ( .A(n2105), .B(n3604), .Z(N10358) );
  CFA1X1 \r347/U1_2  ( .A(n3896), .B(n3771), .CI(\r347/carry [2]), .CO(
        \r347/carry [3]), .S(N6224) );
  CFA1X1 \r347/U1_3  ( .A(n3893), .B(n3270), .CI(\r347/carry [3]), .CO(
        \r347/carry [4]), .S(N6225) );
  CFD2QX1 \lenin0_reg[2]  ( .D(reqlen[2]), .CP(clk), .CD(n3960), .Q(lenin0[2])
         );
  CFD2QXL \wr_ptr_reg[3]  ( .D(N10351), .CP(clk), .CD(n3953), .Q(N2069) );
  CFD2QX1 \wr_ptr_reg[4]  ( .D(N10352), .CP(clk), .CD(n3953), .Q(N2070) );
  CFD2QXL \mem_data1_reg[379]  ( .D(N9703), .CP(clk), .CD(n3962), .Q(
        mem_data1[379]) );
  CFD2QXL \mem_data1_reg[355]  ( .D(N9679), .CP(clk), .CD(n3981), .Q(
        mem_data1[355]) );
  CFD2QXL \mem_data1_reg[357]  ( .D(N9681), .CP(clk), .CD(n3981), .Q(
        mem_data1[357]) );
  CFD2QXL \mem_data1_reg[356]  ( .D(N9680), .CP(clk), .CD(n3981), .Q(
        mem_data1[356]) );
  CFD2QXL \mem_data1_reg[358]  ( .D(N9682), .CP(clk), .CD(n3981), .Q(
        mem_data1[358]) );
  CFD2QXL \mem_data1_reg[352]  ( .D(N9676), .CP(clk), .CD(n3981), .Q(
        mem_data1[352]) );
  CFD2QXL \mem_data1_reg[351]  ( .D(N9675), .CP(clk), .CD(n3980), .Q(
        mem_data1[351]) );
  CFD2QXL \mem_data1_reg[347]  ( .D(N9671), .CP(clk), .CD(n3980), .Q(
        mem_data1[347]) );
  CFD2QXL \mem_data1_reg[380]  ( .D(N9704), .CP(clk), .CD(n3962), .Q(
        mem_data1[380]) );
  CFD2QXL \mem_data1_reg[381]  ( .D(N9705), .CP(clk), .CD(n3962), .Q(
        mem_data1[381]) );
  CFD2QXL \mem_data1_reg[376]  ( .D(N9700), .CP(clk), .CD(n3962), .Q(
        mem_data1[376]) );
  CFD2QXL \mem_data1_reg[413]  ( .D(N9737), .CP(clk), .CD(n3964), .Q(
        mem_data1[413]) );
  CFD2QXL \mem_data1_reg[432]  ( .D(N9756), .CP(clk), .CD(n3966), .Q(
        mem_data1[432]) );
  CFD2QXL \mem_data1_reg[317]  ( .D(N9641), .CP(clk), .CD(n3978), .Q(
        mem_data1[317]) );
  CFD2QXL \mem_data1_reg[315]  ( .D(N9639), .CP(clk), .CD(n3978), .Q(
        mem_data1[315]) );
  CFD2QXL \mem_data1_reg[492]  ( .D(N9816), .CP(clk), .CD(n3971), .Q(
        mem_data1[492]) );
  CFD2QXL \mem_data1_reg[493]  ( .D(N9817), .CP(clk), .CD(n3971), .Q(
        mem_data1[493]) );
  CFD2QXL \mem_data1_reg[491]  ( .D(N9815), .CP(clk), .CD(n3971), .Q(
        mem_data1[491]) );
  CFD2QXL \mem_data1_reg[445]  ( .D(N9769), .CP(clk), .CD(n3967), .Q(
        mem_data1[445]) );
  CFD2QXL \mem_data1_reg[246]  ( .D(N9570), .CP(clk), .CD(n3972), .Q(
        mem_data1[246]) );
  CFD2QXL \mem_data1_reg[290]  ( .D(N9614), .CP(clk), .CD(n3976), .Q(
        mem_data1[290]) );
  CFD2QXL \mem_data1_reg[416]  ( .D(N9740), .CP(clk), .CD(n3965), .Q(
        mem_data1[416]) );
  CFD2QXL \mem_data1_reg[305]  ( .D(N9629), .CP(clk), .CD(n3977), .Q(
        mem_data1[305]) );
  CFD2QXL \mem_data1_reg[303]  ( .D(N9627), .CP(clk), .CD(n3977), .Q(
        mem_data1[303]) );
  CFD2QXL \mem_data1_reg[293]  ( .D(N9617), .CP(clk), .CD(n3976), .Q(
        mem_data1[293]) );
  CFD2QXL \mem_data1_reg[294]  ( .D(N9618), .CP(clk), .CD(n3976), .Q(
        mem_data1[294]) );
  CFD2QXL \mem_data1_reg[292]  ( .D(N9616), .CP(clk), .CD(n3976), .Q(
        mem_data1[292]) );
  CFD2QXL \lenin01_reg[0]  ( .D(n4293), .CP(clk), .CD(n3929), .Q(lenout[0]) );
  CFD2QXL \lenin01_reg[2]  ( .D(n3777), .CP(clk), .CD(n3929), .Q(lenout[2]) );
  CFD2QXL \mem_data1_reg[0]  ( .D(N9324), .CP(clk), .CD(n3953), .Q(
        mem_data1[0]) );
  CFD2QXL \mem_data1_reg[94]  ( .D(N9418), .CP(clk), .CD(n3940), .Q(
        mem_data1[94]) );
  CFD2QXL \mem_data1_reg[102]  ( .D(N9426), .CP(clk), .CD(n3941), .Q(
        mem_data1[102]) );
  CFD2QXL \mem_data1_reg[110]  ( .D(N9434), .CP(clk), .CD(n3941), .Q(
        mem_data1[110]) );
  CFD2QXL \mem_data1_reg[115]  ( .D(N9439), .CP(clk), .CD(n3942), .Q(
        mem_data1[115]) );
  CFD2QXL \mem_data1_reg[116]  ( .D(N9440), .CP(clk), .CD(n3942), .Q(
        mem_data1[116]) );
  CFD2QXL \mem_data1_reg[118]  ( .D(N9442), .CP(clk), .CD(n3942), .Q(
        mem_data1[118]) );
  CFD2QXL \mem_data1_reg[120]  ( .D(N9444), .CP(clk), .CD(n3942), .Q(
        mem_data1[120]) );
  CFD2QXL \mem_data1_reg[230]  ( .D(N9554), .CP(clk), .CD(n3971), .Q(
        mem_data1[230]) );
  CFD2QXL \mem_data1_reg[238]  ( .D(N9562), .CP(clk), .CD(n3972), .Q(
        mem_data1[238]) );
  CFD2QXL \mem_data1_reg[243]  ( .D(N9567), .CP(clk), .CD(n3972), .Q(
        mem_data1[243]) );
  CFD2QXL \mem_data1_reg[245]  ( .D(N9569), .CP(clk), .CD(n3972), .Q(
        mem_data1[245]) );
  CFD2QXL \mem_data1_reg[248]  ( .D(N9572), .CP(clk), .CD(n3973), .Q(
        mem_data1[248]) );
  CFD2QXL \mem_data1_reg[249]  ( .D(N9573), .CP(clk), .CD(n3973), .Q(
        mem_data1[249]) );
  CFD2QXL \mem_data1_reg[250]  ( .D(N9574), .CP(clk), .CD(n3973), .Q(
        mem_data1[250]) );
  CFD2QXL \mem_data1_reg[251]  ( .D(N9575), .CP(clk), .CD(n3973), .Q(
        mem_data1[251]) );
  CFD2QXL \mem_data1_reg[252]  ( .D(N9576), .CP(clk), .CD(n3973), .Q(
        mem_data1[252]) );
  CFD2QXL \mem_data1_reg[353]  ( .D(N9677), .CP(clk), .CD(n3981), .Q(
        mem_data1[353]) );
  CFD2QXL \mem_data1_reg[354]  ( .D(N9678), .CP(clk), .CD(n3981), .Q(
        mem_data1[354]) );
  CFD2QXL \mem_data1_reg[359]  ( .D(N9683), .CP(clk), .CD(n3981), .Q(
        mem_data1[359]) );
  CFD2QXL \mem_data1_reg[361]  ( .D(N9685), .CP(clk), .CD(n3960), .Q(
        mem_data1[361]) );
  CFD2QXL \mem_data1_reg[362]  ( .D(N9686), .CP(clk), .CD(n3961), .Q(
        mem_data1[362]) );
  CFD2QXL \mem_data1_reg[363]  ( .D(N9687), .CP(clk), .CD(n3961), .Q(
        mem_data1[363]) );
  CFD2QXL \mem_data1_reg[366]  ( .D(N9690), .CP(clk), .CD(n3961), .Q(
        mem_data1[366]) );
  CFD2QXL \mem_data1_reg[367]  ( .D(N9691), .CP(clk), .CD(n3961), .Q(
        mem_data1[367]) );
  CFD2QXL \mem_data1_reg[369]  ( .D(N9693), .CP(clk), .CD(n3961), .Q(
        mem_data1[369]) );
  CFD2QXL \mem_data1_reg[373]  ( .D(N9697), .CP(clk), .CD(n3961), .Q(
        mem_data1[373]) );
  CFD2QXL \mem_data1_reg[374]  ( .D(N9698), .CP(clk), .CD(n3961), .Q(
        mem_data1[374]) );
  CFD2QXL \mem_data1_reg[377]  ( .D(N9701), .CP(clk), .CD(n3962), .Q(
        mem_data1[377]) );
  CFD2QXL \mem_data1_reg[483]  ( .D(N9807), .CP(clk), .CD(n3970), .Q(
        mem_data1[483]) );
  CFD2QXL \mem_data1_reg[486]  ( .D(N9810), .CP(clk), .CD(n3970), .Q(
        mem_data1[486]) );
  CFD2QXL \mem_data1_reg[488]  ( .D(N9812), .CP(clk), .CD(n3970), .Q(
        mem_data1[488]) );
  CFD2QXL \mem_data1_reg[489]  ( .D(N9813), .CP(clk), .CD(n3970), .Q(
        mem_data1[489]) );
  CFD2QXL \mem_data1_reg[490]  ( .D(N9814), .CP(clk), .CD(n3970), .Q(
        mem_data1[490]) );
  CFD2QXL \mem_data1_reg[481]  ( .D(N9805), .CP(clk), .CD(n3970), .Q(
        mem_data1[481]) );
  CFD2QXL \mem_data1_reg[484]  ( .D(N9808), .CP(clk), .CD(n3970), .Q(
        mem_data1[484]) );
  CFD2QXL \mem_data1_reg[99]  ( .D(N9423), .CP(clk), .CD(n3940), .Q(
        mem_data1[99]) );
  CFD2QXL \mem_data1_reg[101]  ( .D(N9425), .CP(clk), .CD(n3940), .Q(
        mem_data1[101]) );
  CFD2QXL \mem_data1_reg[103]  ( .D(N9427), .CP(clk), .CD(n3941), .Q(
        mem_data1[103]) );
  CFD2QXL \mem_data1_reg[104]  ( .D(N9428), .CP(clk), .CD(n3941), .Q(
        mem_data1[104]) );
  CFD2QXL \mem_data1_reg[109]  ( .D(N9433), .CP(clk), .CD(n3941), .Q(
        mem_data1[109]) );
  CFD2QXL \mem_data1_reg[114]  ( .D(N9438), .CP(clk), .CD(n3941), .Q(
        mem_data1[114]) );
  CFD2QXL \mem_data1_reg[117]  ( .D(N9441), .CP(clk), .CD(n3942), .Q(
        mem_data1[117]) );
  CFD2QXL \mem_data1_reg[122]  ( .D(N9446), .CP(clk), .CD(n3942), .Q(
        mem_data1[122]) );
  CFD2QXL \mem_data1_reg[125]  ( .D(N9449), .CP(clk), .CD(n3942), .Q(
        mem_data1[125]) );
  CFD2QXL \mem_data1_reg[126]  ( .D(N9450), .CP(clk), .CD(n3942), .Q(
        mem_data1[126]) );
  CFD2QXL \mem_data1_reg[227]  ( .D(N9551), .CP(clk), .CD(n3971), .Q(
        mem_data1[227]) );
  CFD2QXL \mem_data1_reg[232]  ( .D(N9556), .CP(clk), .CD(n3971), .Q(
        mem_data1[232]) );
  CFD2QXL \mem_data1_reg[239]  ( .D(N9563), .CP(clk), .CD(n3972), .Q(
        mem_data1[239]) );
  CFD2QXL \mem_data1_reg[241]  ( .D(N9565), .CP(clk), .CD(n3972), .Q(
        mem_data1[241]) );
  CFD2QXL \mem_data1_reg[244]  ( .D(N9568), .CP(clk), .CD(n3972), .Q(
        mem_data1[244]) );
  CFD2QXL \mem_data1_reg[247]  ( .D(N9571), .CP(clk), .CD(n3972), .Q(
        mem_data1[247]) );
  CFD2QXL \mem_data1_reg[254]  ( .D(N9578), .CP(clk), .CD(n3973), .Q(
        mem_data1[254]) );
  CFD2QXL \mem_data1_reg[360]  ( .D(N9684), .CP(clk), .CD(n3966), .Q(
        mem_data1[360]) );
  CFD2QXL \mem_data1_reg[364]  ( .D(N9688), .CP(clk), .CD(n3961), .Q(
        mem_data1[364]) );
  CFD2QXL \mem_data1_reg[371]  ( .D(N9695), .CP(clk), .CD(n3961), .Q(
        mem_data1[371]) );
  CFD2QXL \mem_data1_reg[372]  ( .D(N9696), .CP(clk), .CD(n3961), .Q(
        mem_data1[372]) );
  CFD2QXL \mem_data1_reg[375]  ( .D(N9699), .CP(clk), .CD(n3962), .Q(
        mem_data1[375]) );
  CFD2QXL \mem_data1_reg[482]  ( .D(N9806), .CP(clk), .CD(n3970), .Q(
        mem_data1[482]) );
  CFD2QXL \mem_data1_reg[495]  ( .D(N9819), .CP(clk), .CD(n3919), .Q(
        mem_data1[495]) );
  CFD2QXL \mem_data1_reg[496]  ( .D(N9820), .CP(clk), .CD(n3914), .Q(
        mem_data1[496]) );
  CFD2QXL \mem_data1_reg[499]  ( .D(N9823), .CP(clk), .CD(n3909), .Q(
        mem_data1[499]) );
  CFD2QXL \mem_data1_reg[33]  ( .D(N9357), .CP(clk), .CD(n3956), .Q(
        mem_data1[33]) );
  CFD2QXL \mem_data1_reg[58]  ( .D(N9382), .CP(clk), .CD(n3958), .Q(
        mem_data1[58]) );
  CFD2QXL \mem_data1_reg[59]  ( .D(N9383), .CP(clk), .CD(n3958), .Q(
        mem_data1[59]) );
  CFD2QXL \mem_data1_reg[61]  ( .D(N9385), .CP(clk), .CD(n3958), .Q(
        mem_data1[61]) );
  CFD2QXL \mem_data1_reg[90]  ( .D(N9414), .CP(clk), .CD(n3945), .Q(
        mem_data1[90]) );
  CFD2QXL \mem_data1_reg[98]  ( .D(N9422), .CP(clk), .CD(n3940), .Q(
        mem_data1[98]) );
  CFD2QXL \mem_data1_reg[111]  ( .D(N9435), .CP(clk), .CD(n3941), .Q(
        mem_data1[111]) );
  CFD2QXL \mem_data1_reg[112]  ( .D(N9436), .CP(clk), .CD(n3941), .Q(
        mem_data1[112]) );
  CFD2QXL \mem_data1_reg[113]  ( .D(N9437), .CP(clk), .CD(n3941), .Q(
        mem_data1[113]) );
  CFD2QXL \mem_data1_reg[119]  ( .D(N9443), .CP(clk), .CD(n3942), .Q(
        mem_data1[119]) );
  CFD2QXL \mem_data1_reg[123]  ( .D(N9447), .CP(clk), .CD(n3942), .Q(
        mem_data1[123]) );
  CFD2QXL \mem_data1_reg[156]  ( .D(N9480), .CP(clk), .CD(n3945), .Q(
        mem_data1[156]) );
  CFD2QXL \mem_data1_reg[162]  ( .D(N9486), .CP(clk), .CD(n3945), .Q(
        mem_data1[162]) );
  CFD2QXL \mem_data1_reg[181]  ( .D(N9505), .CP(clk), .CD(n3947), .Q(
        mem_data1[181]) );
  CFD2QXL \mem_data1_reg[182]  ( .D(N9506), .CP(clk), .CD(n3947), .Q(
        mem_data1[182]) );
  CFD2QXL \mem_data1_reg[183]  ( .D(N9507), .CP(clk), .CD(n3947), .Q(
        mem_data1[183]) );
  CFD2QXL \mem_data1_reg[185]  ( .D(N9509), .CP(clk), .CD(n3947), .Q(
        mem_data1[185]) );
  CFD2QXL \mem_data1_reg[186]  ( .D(N9510), .CP(clk), .CD(n3947), .Q(
        mem_data1[186]) );
  CFD2QXL \mem_data1_reg[187]  ( .D(N9511), .CP(clk), .CD(n3947), .Q(
        mem_data1[187]) );
  CFD2QXL \mem_data1_reg[189]  ( .D(N9513), .CP(clk), .CD(n3947), .Q(
        mem_data1[189]) );
  CFD2QXL \mem_data1_reg[220]  ( .D(N9544), .CP(clk), .CD(n3950), .Q(
        mem_data1[220]) );
  CFD2QXL \mem_data1_reg[228]  ( .D(N9552), .CP(clk), .CD(n3971), .Q(
        mem_data1[228]) );
  CFD2QXL \mem_data1_reg[234]  ( .D(N9558), .CP(clk), .CD(n3971), .Q(
        mem_data1[234]) );
  CFD2QXL \mem_data1_reg[242]  ( .D(N9566), .CP(clk), .CD(n3972), .Q(
        mem_data1[242]) );
  CFD2QXL \mem_data1_reg[256]  ( .D(N9580), .CP(clk), .CD(n3973), .Q(
        mem_data1[256]) );
  CFD2QXL \mem_data1_reg[257]  ( .D(N9581), .CP(clk), .CD(n3973), .Q(
        mem_data1[257]) );
  CFD2QXL \mem_data1_reg[259]  ( .D(N9583), .CP(clk), .CD(n3973), .Q(
        mem_data1[259]) );
  CFD2QXL \mem_data1_reg[261]  ( .D(N9585), .CP(clk), .CD(n3974), .Q(
        mem_data1[261]) );
  CFD2QXL \mem_data1_reg[271]  ( .D(N9595), .CP(clk), .CD(n3974), .Q(
        mem_data1[271]) );
  CFD2QXL \mem_data1_reg[273]  ( .D(N9597), .CP(clk), .CD(n3974), .Q(
        mem_data1[273]) );
  CFD2QXL \mem_data1_reg[277]  ( .D(N9601), .CP(clk), .CD(n3975), .Q(
        mem_data1[277]) );
  CFD2QXL \mem_data1_reg[278]  ( .D(N9602), .CP(clk), .CD(n3975), .Q(
        mem_data1[278]) );
  CFD2QXL \mem_data1_reg[279]  ( .D(N9603), .CP(clk), .CD(n3975), .Q(
        mem_data1[279]) );
  CFD2QXL \mem_data1_reg[282]  ( .D(N9606), .CP(clk), .CD(n3975), .Q(
        mem_data1[282]) );
  CFD2QXL \mem_data1_reg[283]  ( .D(N9607), .CP(clk), .CD(n3975), .Q(
        mem_data1[283]) );
  CFD2QXL \mem_data1_reg[286]  ( .D(N9610), .CP(clk), .CD(n3975), .Q(
        mem_data1[286]) );
  CFD2QXL \mem_data1_reg[299]  ( .D(N9623), .CP(clk), .CD(n3977), .Q(
        mem_data1[299]) );
  CFD2QXL \mem_data1_reg[301]  ( .D(N9625), .CP(clk), .CD(n3977), .Q(
        mem_data1[301]) );
  CFD2QXL \mem_data1_reg[304]  ( .D(N9628), .CP(clk), .CD(n3977), .Q(
        mem_data1[304]) );
  CFD2QXL \mem_data1_reg[309]  ( .D(N9633), .CP(clk), .CD(n3977), .Q(
        mem_data1[309]) );
  CFD2QXL \mem_data1_reg[313]  ( .D(N9637), .CP(clk), .CD(n3978), .Q(
        mem_data1[313]) );
  CFD2QXL \mem_data1_reg[314]  ( .D(N9638), .CP(clk), .CD(n3978), .Q(
        mem_data1[314]) );
  CFD2QXL \mem_data1_reg[316]  ( .D(N9640), .CP(clk), .CD(n3978), .Q(
        mem_data1[316]) );
  CFD2QXL \mem_data1_reg[320]  ( .D(N9644), .CP(clk), .CD(n3978), .Q(
        mem_data1[320]) );
  CFD2QXL \mem_data1_reg[321]  ( .D(N9645), .CP(clk), .CD(n3978), .Q(
        mem_data1[321]) );
  CFD2QXL \mem_data1_reg[323]  ( .D(N9647), .CP(clk), .CD(n3978), .Q(
        mem_data1[323]) );
  CFD2QXL \mem_data1_reg[324]  ( .D(N9648), .CP(clk), .CD(n3979), .Q(
        mem_data1[324]) );
  CFD2QXL \mem_data1_reg[325]  ( .D(N9649), .CP(clk), .CD(n3978), .Q(
        mem_data1[325]) );
  CFD2QXL \mem_data1_reg[326]  ( .D(N9650), .CP(clk), .CD(n3979), .Q(
        mem_data1[326]) );
  CFD2QXL \mem_data1_reg[327]  ( .D(N9651), .CP(clk), .CD(n3979), .Q(
        mem_data1[327]) );
  CFD2QXL \mem_data1_reg[335]  ( .D(N9659), .CP(clk), .CD(n3979), .Q(
        mem_data1[335]) );
  CFD2QXL \mem_data1_reg[339]  ( .D(N9663), .CP(clk), .CD(n3979), .Q(
        mem_data1[339]) );
  CFD2QXL \mem_data1_reg[340]  ( .D(N9664), .CP(clk), .CD(n3980), .Q(
        mem_data1[340]) );
  CFD2QXL \mem_data1_reg[341]  ( .D(N9665), .CP(clk), .CD(n3980), .Q(
        mem_data1[341]) );
  CFD2QXL \mem_data1_reg[342]  ( .D(N9666), .CP(clk), .CD(n3980), .Q(
        mem_data1[342]) );
  CFD2QXL \mem_data1_reg[343]  ( .D(N9667), .CP(clk), .CD(n3980), .Q(
        mem_data1[343]) );
  CFD2QXL \mem_data1_reg[344]  ( .D(N9668), .CP(clk), .CD(n3980), .Q(
        mem_data1[344]) );
  CFD2QXL \mem_data1_reg[345]  ( .D(N9669), .CP(clk), .CD(n3980), .Q(
        mem_data1[345]) );
  CFD2QXL \mem_data1_reg[346]  ( .D(N9670), .CP(clk), .CD(n3980), .Q(
        mem_data1[346]) );
  CFD2QXL \mem_data1_reg[348]  ( .D(N9672), .CP(clk), .CD(n3980), .Q(
        mem_data1[348]) );
  CFD2QXL \mem_data1_reg[349]  ( .D(N9673), .CP(clk), .CD(n3980), .Q(
        mem_data1[349]) );
  CFD2QXL \mem_data1_reg[350]  ( .D(N9674), .CP(clk), .CD(n3981), .Q(
        mem_data1[350]) );
  CFD2QXL \mem_data1_reg[365]  ( .D(N9689), .CP(clk), .CD(n3961), .Q(
        mem_data1[365]) );
  CFD2QXL \mem_data1_reg[370]  ( .D(N9694), .CP(clk), .CD(n3961), .Q(
        mem_data1[370]) );
  CFD2QXL \mem_data1_reg[378]  ( .D(N9702), .CP(clk), .CD(n3962), .Q(
        mem_data1[378]) );
  CFD2QXL \mem_data1_reg[385]  ( .D(N9709), .CP(clk), .CD(n3962), .Q(
        mem_data1[385]) );
  CFD2QXL \mem_data1_reg[386]  ( .D(N9710), .CP(clk), .CD(n3962), .Q(
        mem_data1[386]) );
  CFD2QXL \mem_data1_reg[387]  ( .D(N9711), .CP(clk), .CD(n3962), .Q(
        mem_data1[387]) );
  CFD2QXL \mem_data1_reg[388]  ( .D(N9712), .CP(clk), .CD(n3963), .Q(
        mem_data1[388]) );
  CFD2QXL \mem_data1_reg[389]  ( .D(N9713), .CP(clk), .CD(n3963), .Q(
        mem_data1[389]) );
  CFD2QXL \mem_data1_reg[391]  ( .D(N9715), .CP(clk), .CD(n3963), .Q(
        mem_data1[391]) );
  CFD2QXL \mem_data1_reg[393]  ( .D(N9717), .CP(clk), .CD(n3963), .Q(
        mem_data1[393]) );
  CFD2QXL \mem_data1_reg[395]  ( .D(N9719), .CP(clk), .CD(n3963), .Q(
        mem_data1[395]) );
  CFD2QXL \mem_data1_reg[396]  ( .D(N9720), .CP(clk), .CD(n3963), .Q(
        mem_data1[396]) );
  CFD2QXL \mem_data1_reg[397]  ( .D(N9721), .CP(clk), .CD(n3963), .Q(
        mem_data1[397]) );
  CFD2QXL \mem_data1_reg[398]  ( .D(N9722), .CP(clk), .CD(n3963), .Q(
        mem_data1[398]) );
  CFD2QXL \mem_data1_reg[399]  ( .D(N9723), .CP(clk), .CD(n3963), .Q(
        mem_data1[399]) );
  CFD2QXL \mem_data1_reg[401]  ( .D(N9725), .CP(clk), .CD(n3964), .Q(
        mem_data1[401]) );
  CFD2QXL \mem_data1_reg[402]  ( .D(N9726), .CP(clk), .CD(n3964), .Q(
        mem_data1[402]) );
  CFD2QXL \mem_data1_reg[404]  ( .D(N9728), .CP(clk), .CD(n3964), .Q(
        mem_data1[404]) );
  CFD2QXL \mem_data1_reg[405]  ( .D(N9729), .CP(clk), .CD(n3964), .Q(
        mem_data1[405]) );
  CFD2QXL \mem_data1_reg[407]  ( .D(N9731), .CP(clk), .CD(n3964), .Q(
        mem_data1[407]) );
  CFD2QXL \mem_data1_reg[408]  ( .D(N9732), .CP(clk), .CD(n3964), .Q(
        mem_data1[408]) );
  CFD2QXL \mem_data1_reg[409]  ( .D(N9733), .CP(clk), .CD(n3964), .Q(
        mem_data1[409]) );
  CFD2QXL \mem_data1_reg[410]  ( .D(N9734), .CP(clk), .CD(n3964), .Q(
        mem_data1[410]) );
  CFD2QXL \mem_data1_reg[411]  ( .D(N9735), .CP(clk), .CD(n3964), .Q(
        mem_data1[411]) );
  CFD2QXL \mem_data1_reg[412]  ( .D(N9736), .CP(clk), .CD(n3964), .Q(
        mem_data1[412]) );
  CFD2QXL \mem_data1_reg[415]  ( .D(N9739), .CP(clk), .CD(n3965), .Q(
        mem_data1[415]) );
  CFD2QXL \mem_data1_reg[425]  ( .D(N9749), .CP(clk), .CD(n3965), .Q(
        mem_data1[425]) );
  CFD2QXL \mem_data1_reg[426]  ( .D(N9750), .CP(clk), .CD(n3965), .Q(
        mem_data1[426]) );
  CFD2QXL \mem_data1_reg[428]  ( .D(N9752), .CP(clk), .CD(n3966), .Q(
        mem_data1[428]) );
  CFD2QXL \mem_data1_reg[429]  ( .D(N9753), .CP(clk), .CD(n3966), .Q(
        mem_data1[429]) );
  CFD2QXL \mem_data1_reg[434]  ( .D(N9758), .CP(clk), .CD(n3966), .Q(
        mem_data1[434]) );
  CFD2QXL \mem_data1_reg[438]  ( .D(N9762), .CP(clk), .CD(n3966), .Q(
        mem_data1[438]) );
  CFD2QXL \mem_data1_reg[439]  ( .D(N9763), .CP(clk), .CD(n3967), .Q(
        mem_data1[439]) );
  CFD2QXL \mem_data1_reg[440]  ( .D(N9764), .CP(clk), .CD(n3967), .Q(
        mem_data1[440]) );
  CFD2QXL \mem_data1_reg[450]  ( .D(N9774), .CP(clk), .CD(n3967), .Q(
        mem_data1[450]) );
  CFD2QXL \mem_data1_reg[451]  ( .D(N9775), .CP(clk), .CD(n3967), .Q(
        mem_data1[451]) );
  CFD2QXL \mem_data1_reg[453]  ( .D(N9777), .CP(clk), .CD(n3968), .Q(
        mem_data1[453]) );
  CFD2QXL \mem_data1_reg[455]  ( .D(N9779), .CP(clk), .CD(n3968), .Q(
        mem_data1[455]) );
  CFD2QXL \mem_data1_reg[457]  ( .D(N9781), .CP(clk), .CD(n3968), .Q(
        mem_data1[457]) );
  CFD2QXL \mem_data1_reg[460]  ( .D(N9784), .CP(clk), .CD(n3968), .Q(
        mem_data1[460]) );
  CFD2QXL \mem_data1_reg[461]  ( .D(N9785), .CP(clk), .CD(n3968), .Q(
        mem_data1[461]) );
  CFD2QXL \mem_data1_reg[463]  ( .D(N9787), .CP(clk), .CD(n3968), .Q(
        mem_data1[463]) );
  CFD2QXL \mem_data1_reg[464]  ( .D(N9788), .CP(clk), .CD(n3968), .Q(
        mem_data1[464]) );
  CFD2QXL \mem_data1_reg[465]  ( .D(N9789), .CP(clk), .CD(n3969), .Q(
        mem_data1[465]) );
  CFD2QXL \mem_data1_reg[469]  ( .D(N9793), .CP(clk), .CD(n3969), .Q(
        mem_data1[469]) );
  CFD2QXL \mem_data1_reg[473]  ( .D(N9797), .CP(clk), .CD(n3969), .Q(
        mem_data1[473]) );
  CFD2QXL \mem_data1_reg[475]  ( .D(N9799), .CP(clk), .CD(n3969), .Q(
        mem_data1[475]) );
  CFD2QXL \mem_data1_reg[477]  ( .D(N9801), .CP(clk), .CD(n3969), .Q(
        mem_data1[477]) );
  CFD2QXL \mem_data1_reg[480]  ( .D(N9804), .CP(clk), .CD(n3970), .Q(
        mem_data1[480]) );
  CFD2QXL \mem_data1_reg[957]  ( .D(N10281), .CP(clk), .CD(n3924), .Q(
        mem_data1[957]) );
  CFD2QXL \mem_data1_reg[295]  ( .D(N9619), .CP(clk), .CD(n3976), .Q(
        mem_data1[295]) );
  CFD2QXL \mem_data1_reg[296]  ( .D(N9620), .CP(clk), .CD(n3976), .Q(
        mem_data1[296]) );
  CFD2QXL \mem_data1_reg[337]  ( .D(N9661), .CP(clk), .CD(n3979), .Q(
        mem_data1[337]) );
  CFD2QXL \mem_data1_reg[421]  ( .D(N9745), .CP(clk), .CD(n3965), .Q(
        mem_data1[421]) );
  CFD2QXL \mem_data1_reg[423]  ( .D(N9747), .CP(clk), .CD(n3965), .Q(
        mem_data1[423]) );
  CFD2QXL \mem_data1_reg[427]  ( .D(N9751), .CP(clk), .CD(n3966), .Q(
        mem_data1[427]) );
  CFD2QXL \mem_data1_reg[430]  ( .D(N9754), .CP(clk), .CD(n3966), .Q(
        mem_data1[430]) );
  CFD2QXL \mem_data1_reg[431]  ( .D(N9755), .CP(clk), .CD(n3966), .Q(
        mem_data1[431]) );
  CFD2QXL \mem_data1_reg[433]  ( .D(N9757), .CP(clk), .CD(n3966), .Q(
        mem_data1[433]) );
  CFD2QXL \mem_data1_reg[435]  ( .D(N9759), .CP(clk), .CD(n3966), .Q(
        mem_data1[435]) );
  CFD2QXL \mem_data1_reg[1023]  ( .D(N10347), .CP(clk), .CD(n3953), .Q(
        mem_data1[1023]) );
  CFD2QXL \mem_data1_reg[676]  ( .D(N10000), .CP(clk), .CD(n3953), .Q(
        mem_data1[676]) );
  CFD2QXL \mem_data1_reg[1022]  ( .D(N10346), .CP(clk), .CD(n3953), .Q(
        mem_data1[1022]) );
  CFD2QXL \mem_data1_reg[15]  ( .D(N9339), .CP(clk), .CD(n3955), .Q(
        mem_data1[15]) );
  CFD2QXL \mem_data1_reg[16]  ( .D(N9340), .CP(clk), .CD(n3955), .Q(
        mem_data1[16]) );
  CFD2QXL \mem_data1_reg[17]  ( .D(N9341), .CP(clk), .CD(n3955), .Q(
        mem_data1[17]) );
  CFD2QXL \mem_data1_reg[18]  ( .D(N9342), .CP(clk), .CD(n3955), .Q(
        mem_data1[18]) );
  CFD2QXL \mem_data1_reg[19]  ( .D(N9343), .CP(clk), .CD(n3955), .Q(
        mem_data1[19]) );
  CFD2QXL \mem_data1_reg[20]  ( .D(N9344), .CP(clk), .CD(n3955), .Q(
        mem_data1[20]) );
  CFD2QXL \mem_data1_reg[21]  ( .D(N9345), .CP(clk), .CD(n3955), .Q(
        mem_data1[21]) );
  CFD2QXL \mem_data1_reg[22]  ( .D(N9346), .CP(clk), .CD(n3955), .Q(
        mem_data1[22]) );
  CFD2QXL \mem_data1_reg[23]  ( .D(N9347), .CP(clk), .CD(n3955), .Q(
        mem_data1[23]) );
  CFD2QXL \mem_data1_reg[24]  ( .D(N9348), .CP(clk), .CD(n3955), .Q(
        mem_data1[24]) );
  CFD2QXL \mem_data1_reg[25]  ( .D(N9349), .CP(clk), .CD(n3955), .Q(
        mem_data1[25]) );
  CFD2QXL \mem_data1_reg[26]  ( .D(N9350), .CP(clk), .CD(n3955), .Q(
        mem_data1[26]) );
  CFD2QXL \mem_data1_reg[27]  ( .D(N9351), .CP(clk), .CD(n3956), .Q(
        mem_data1[27]) );
  CFD2QXL \mem_data1_reg[28]  ( .D(N9352), .CP(clk), .CD(n3956), .Q(
        mem_data1[28]) );
  CFD2QXL \mem_data1_reg[29]  ( .D(N9353), .CP(clk), .CD(n3956), .Q(
        mem_data1[29]) );
  CFD2QXL \mem_data1_reg[30]  ( .D(N9354), .CP(clk), .CD(n3956), .Q(
        mem_data1[30]) );
  CFD2QXL \mem_data1_reg[31]  ( .D(N9355), .CP(clk), .CD(n3956), .Q(
        mem_data1[31]) );
  CFD2QXL \mem_data1_reg[32]  ( .D(N9356), .CP(clk), .CD(n3956), .Q(
        mem_data1[32]) );
  CFD2QXL \mem_data1_reg[34]  ( .D(N9358), .CP(clk), .CD(n3956), .Q(
        mem_data1[34]) );
  CFD2QXL \mem_data1_reg[35]  ( .D(N9359), .CP(clk), .CD(n3956), .Q(
        mem_data1[35]) );
  CFD2QXL \mem_data1_reg[36]  ( .D(N9360), .CP(clk), .CD(n3956), .Q(
        mem_data1[36]) );
  CFD2QXL \mem_data1_reg[37]  ( .D(N9361), .CP(clk), .CD(n3956), .Q(
        mem_data1[37]) );
  CFD2QXL \mem_data1_reg[38]  ( .D(N9362), .CP(clk), .CD(n3956), .Q(
        mem_data1[38]) );
  CFD2QXL \mem_data1_reg[39]  ( .D(N9363), .CP(clk), .CD(n3956), .Q(
        mem_data1[39]) );
  CFD2QXL \mem_data1_reg[40]  ( .D(N9364), .CP(clk), .CD(n3957), .Q(
        mem_data1[40]) );
  CFD2QXL \mem_data1_reg[41]  ( .D(N9365), .CP(clk), .CD(n3957), .Q(
        mem_data1[41]) );
  CFD2QXL \mem_data1_reg[42]  ( .D(N9366), .CP(clk), .CD(n3957), .Q(
        mem_data1[42]) );
  CFD2QXL \mem_data1_reg[43]  ( .D(N9367), .CP(clk), .CD(n3957), .Q(
        mem_data1[43]) );
  CFD2QXL \mem_data1_reg[44]  ( .D(N9368), .CP(clk), .CD(n3957), .Q(
        mem_data1[44]) );
  CFD2QXL \mem_data1_reg[45]  ( .D(N9369), .CP(clk), .CD(n3957), .Q(
        mem_data1[45]) );
  CFD2QXL \mem_data1_reg[46]  ( .D(N9370), .CP(clk), .CD(n3957), .Q(
        mem_data1[46]) );
  CFD2QXL \mem_data1_reg[47]  ( .D(N9371), .CP(clk), .CD(n3957), .Q(
        mem_data1[47]) );
  CFD2QXL \mem_data1_reg[48]  ( .D(N9372), .CP(clk), .CD(n3957), .Q(
        mem_data1[48]) );
  CFD2QXL \mem_data1_reg[49]  ( .D(N9373), .CP(clk), .CD(n3957), .Q(
        mem_data1[49]) );
  CFD2QXL \mem_data1_reg[50]  ( .D(N9374), .CP(clk), .CD(n3957), .Q(
        mem_data1[50]) );
  CFD2QXL \mem_data1_reg[51]  ( .D(N9375), .CP(clk), .CD(n3957), .Q(
        mem_data1[51]) );
  CFD2QXL \mem_data1_reg[52]  ( .D(N9376), .CP(clk), .CD(n3957), .Q(
        mem_data1[52]) );
  CFD2QXL \mem_data1_reg[53]  ( .D(N9377), .CP(clk), .CD(n3958), .Q(
        mem_data1[53]) );
  CFD2QXL \mem_data1_reg[54]  ( .D(N9378), .CP(clk), .CD(n3958), .Q(
        mem_data1[54]) );
  CFD2QXL \mem_data1_reg[55]  ( .D(N9379), .CP(clk), .CD(n3958), .Q(
        mem_data1[55]) );
  CFD2QXL \mem_data1_reg[56]  ( .D(N9380), .CP(clk), .CD(n3958), .Q(
        mem_data1[56]) );
  CFD2QXL \mem_data1_reg[57]  ( .D(N9381), .CP(clk), .CD(n3958), .Q(
        mem_data1[57]) );
  CFD2QXL \mem_data1_reg[60]  ( .D(N9384), .CP(clk), .CD(n3958), .Q(
        mem_data1[60]) );
  CFD2QXL \mem_data1_reg[62]  ( .D(N9386), .CP(clk), .CD(n3958), .Q(
        mem_data1[62]) );
  CFD2QXL \mem_data1_reg[63]  ( .D(N9387), .CP(clk), .CD(n3958), .Q(
        mem_data1[63]) );
  CFD2QXL \mem_data1_reg[64]  ( .D(N9388), .CP(clk), .CD(n3958), .Q(
        mem_data1[64]) );
  CFD2QXL \mem_data1_reg[65]  ( .D(N9389), .CP(clk), .CD(n3958), .Q(
        mem_data1[65]) );
  CFD2QXL \mem_data1_reg[66]  ( .D(N9390), .CP(clk), .CD(n3959), .Q(
        mem_data1[66]) );
  CFD2QXL \mem_data1_reg[67]  ( .D(N9391), .CP(clk), .CD(n3959), .Q(
        mem_data1[67]) );
  CFD2QXL \mem_data1_reg[68]  ( .D(N9392), .CP(clk), .CD(n3959), .Q(
        mem_data1[68]) );
  CFD2QXL \mem_data1_reg[69]  ( .D(N9393), .CP(clk), .CD(n3959), .Q(
        mem_data1[69]) );
  CFD2QXL \mem_data1_reg[70]  ( .D(N9394), .CP(clk), .CD(n3959), .Q(
        mem_data1[70]) );
  CFD2QXL \mem_data1_reg[71]  ( .D(N9395), .CP(clk), .CD(n3959), .Q(
        mem_data1[71]) );
  CFD2QXL \mem_data1_reg[72]  ( .D(N9396), .CP(clk), .CD(n3959), .Q(
        mem_data1[72]) );
  CFD2QXL \mem_data1_reg[73]  ( .D(N9397), .CP(clk), .CD(n3959), .Q(
        mem_data1[73]) );
  CFD2QXL \mem_data1_reg[74]  ( .D(N9398), .CP(clk), .CD(n3959), .Q(
        mem_data1[74]) );
  CFD2QXL \mem_data1_reg[75]  ( .D(N9399), .CP(clk), .CD(n3959), .Q(
        mem_data1[75]) );
  CFD2QXL \mem_data1_reg[76]  ( .D(N9400), .CP(clk), .CD(n3959), .Q(
        mem_data1[76]) );
  CFD2QXL \mem_data1_reg[77]  ( .D(N9401), .CP(clk), .CD(n3959), .Q(
        mem_data1[77]) );
  CFD2QXL \mem_data1_reg[78]  ( .D(N9402), .CP(clk), .CD(n3959), .Q(
        mem_data1[78]) );
  CFD2QXL \mem_data1_reg[79]  ( .D(N9403), .CP(clk), .CD(n3960), .Q(
        mem_data1[79]) );
  CFD2QXL \mem_data1_reg[80]  ( .D(N9404), .CP(clk), .CD(n3960), .Q(
        mem_data1[80]) );
  CFD2QXL \mem_data1_reg[81]  ( .D(N9405), .CP(clk), .CD(n3960), .Q(
        mem_data1[81]) );
  CFD2QXL \mem_data1_reg[82]  ( .D(N9406), .CP(clk), .CD(n3960), .Q(
        mem_data1[82]) );
  CFD2QXL \mem_data1_reg[83]  ( .D(N9407), .CP(clk), .CD(n3960), .Q(
        mem_data1[83]) );
  CFD2QXL \mem_data1_reg[84]  ( .D(N9408), .CP(clk), .CD(n3960), .Q(
        mem_data1[84]) );
  CFD2QXL \mem_data1_reg[85]  ( .D(N9409), .CP(clk), .CD(n3960), .Q(
        mem_data1[85]) );
  CFD2QXL \mem_data1_reg[86]  ( .D(N9410), .CP(clk), .CD(n3960), .Q(
        mem_data1[86]) );
  CFD2QXL \mem_data1_reg[87]  ( .D(N9411), .CP(clk), .CD(n3960), .Q(
        mem_data1[87]) );
  CFD2QXL \mem_data1_reg[88]  ( .D(N9412), .CP(clk), .CD(n3960), .Q(
        mem_data1[88]) );
  CFD2QXL \mem_data1_reg[89]  ( .D(N9413), .CP(clk), .CD(n3960), .Q(
        mem_data1[89]) );
  CFD2QXL \mem_data1_reg[91]  ( .D(N9415), .CP(clk), .CD(n3940), .Q(
        mem_data1[91]) );
  CFD2QXL \mem_data1_reg[92]  ( .D(N9416), .CP(clk), .CD(n3940), .Q(
        mem_data1[92]) );
  CFD2QXL \mem_data1_reg[93]  ( .D(N9417), .CP(clk), .CD(n3940), .Q(
        mem_data1[93]) );
  CFD2QXL \mem_data1_reg[95]  ( .D(N9419), .CP(clk), .CD(n3940), .Q(
        mem_data1[95]) );
  CFD2QXL \mem_data1_reg[96]  ( .D(N9420), .CP(clk), .CD(n3940), .Q(
        mem_data1[96]) );
  CFD2QXL \mem_data1_reg[97]  ( .D(N9421), .CP(clk), .CD(n3940), .Q(
        mem_data1[97]) );
  CFD2QXL \mem_data1_reg[100]  ( .D(N9424), .CP(clk), .CD(n3940), .Q(
        mem_data1[100]) );
  CFD2QXL \mem_data1_reg[105]  ( .D(N9429), .CP(clk), .CD(n3941), .Q(
        mem_data1[105]) );
  CFD2QXL \mem_data1_reg[106]  ( .D(N9430), .CP(clk), .CD(n3941), .Q(
        mem_data1[106]) );
  CFD2QXL \mem_data1_reg[107]  ( .D(N9431), .CP(clk), .CD(n3941), .Q(
        mem_data1[107]) );
  CFD2QXL \mem_data1_reg[108]  ( .D(N9432), .CP(clk), .CD(n3941), .Q(
        mem_data1[108]) );
  CFD2QXL \mem_data1_reg[121]  ( .D(N9445), .CP(clk), .CD(n3942), .Q(
        mem_data1[121]) );
  CFD2QXL \mem_data1_reg[124]  ( .D(N9448), .CP(clk), .CD(n3942), .Q(
        mem_data1[124]) );
  CFD2QXL \mem_data1_reg[127]  ( .D(N9451), .CP(clk), .CD(n3942), .Q(
        mem_data1[127]) );
  CFD2QXL \mem_data1_reg[128]  ( .D(N9452), .CP(clk), .CD(n3943), .Q(
        mem_data1[128]) );
  CFD2QXL \mem_data1_reg[129]  ( .D(N9453), .CP(clk), .CD(n3943), .Q(
        mem_data1[129]) );
  CFD2QXL \mem_data1_reg[130]  ( .D(N9454), .CP(clk), .CD(n3943), .Q(
        mem_data1[130]) );
  CFD2QXL \mem_data1_reg[131]  ( .D(N9455), .CP(clk), .CD(n3943), .Q(
        mem_data1[131]) );
  CFD2QXL \mem_data1_reg[132]  ( .D(N9456), .CP(clk), .CD(n3943), .Q(
        mem_data1[132]) );
  CFD2QXL \mem_data1_reg[133]  ( .D(N9457), .CP(clk), .CD(n3943), .Q(
        mem_data1[133]) );
  CFD2QXL \mem_data1_reg[134]  ( .D(N9458), .CP(clk), .CD(n3943), .Q(
        mem_data1[134]) );
  CFD2QXL \mem_data1_reg[135]  ( .D(N9459), .CP(clk), .CD(n3943), .Q(
        mem_data1[135]) );
  CFD2QXL \mem_data1_reg[136]  ( .D(N9460), .CP(clk), .CD(n3943), .Q(
        mem_data1[136]) );
  CFD2QXL \mem_data1_reg[137]  ( .D(N9461), .CP(clk), .CD(n3943), .Q(
        mem_data1[137]) );
  CFD2QXL \mem_data1_reg[138]  ( .D(N9462), .CP(clk), .CD(n3943), .Q(
        mem_data1[138]) );
  CFD2QXL \mem_data1_reg[139]  ( .D(N9463), .CP(clk), .CD(n3943), .Q(
        mem_data1[139]) );
  CFD2QXL \mem_data1_reg[140]  ( .D(N9464), .CP(clk), .CD(n3943), .Q(
        mem_data1[140]) );
  CFD2QXL \mem_data1_reg[141]  ( .D(N9465), .CP(clk), .CD(n3944), .Q(
        mem_data1[141]) );
  CFD2QXL \mem_data1_reg[142]  ( .D(N9466), .CP(clk), .CD(n3944), .Q(
        mem_data1[142]) );
  CFD2QXL \mem_data1_reg[143]  ( .D(N9467), .CP(clk), .CD(n3944), .Q(
        mem_data1[143]) );
  CFD2QXL \mem_data1_reg[144]  ( .D(N9468), .CP(clk), .CD(n3944), .Q(
        mem_data1[144]) );
  CFD2QXL \mem_data1_reg[145]  ( .D(N9469), .CP(clk), .CD(n3944), .Q(
        mem_data1[145]) );
  CFD2QXL \mem_data1_reg[146]  ( .D(N9470), .CP(clk), .CD(n3944), .Q(
        mem_data1[146]) );
  CFD2QXL \mem_data1_reg[147]  ( .D(N9471), .CP(clk), .CD(n3944), .Q(
        mem_data1[147]) );
  CFD2QXL \mem_data1_reg[148]  ( .D(N9472), .CP(clk), .CD(n3944), .Q(
        mem_data1[148]) );
  CFD2QXL \mem_data1_reg[149]  ( .D(N9473), .CP(clk), .CD(n3944), .Q(
        mem_data1[149]) );
  CFD2QXL \mem_data1_reg[150]  ( .D(N9474), .CP(clk), .CD(n3944), .Q(
        mem_data1[150]) );
  CFD2QXL \mem_data1_reg[151]  ( .D(N9475), .CP(clk), .CD(n3944), .Q(
        mem_data1[151]) );
  CFD2QXL \mem_data1_reg[152]  ( .D(N9476), .CP(clk), .CD(n3944), .Q(
        mem_data1[152]) );
  CFD2QXL \mem_data1_reg[153]  ( .D(N9477), .CP(clk), .CD(n3944), .Q(
        mem_data1[153]) );
  CFD2QXL \mem_data1_reg[154]  ( .D(N9478), .CP(clk), .CD(n3945), .Q(
        mem_data1[154]) );
  CFD2QXL \mem_data1_reg[155]  ( .D(N9479), .CP(clk), .CD(n3945), .Q(
        mem_data1[155]) );
  CFD2QXL \mem_data1_reg[157]  ( .D(N9481), .CP(clk), .CD(n3945), .Q(
        mem_data1[157]) );
  CFD2QXL \mem_data1_reg[158]  ( .D(N9482), .CP(clk), .CD(n3945), .Q(
        mem_data1[158]) );
  CFD2QXL \mem_data1_reg[159]  ( .D(N9483), .CP(clk), .CD(n3945), .Q(
        mem_data1[159]) );
  CFD2QXL \mem_data1_reg[160]  ( .D(N9484), .CP(clk), .CD(n3945), .Q(
        mem_data1[160]) );
  CFD2QXL \mem_data1_reg[161]  ( .D(N9485), .CP(clk), .CD(n3945), .Q(
        mem_data1[161]) );
  CFD2QXL \mem_data1_reg[163]  ( .D(N9487), .CP(clk), .CD(n3945), .Q(
        mem_data1[163]) );
  CFD2QXL \mem_data1_reg[164]  ( .D(N9488), .CP(clk), .CD(n3945), .Q(
        mem_data1[164]) );
  CFD2QXL \mem_data1_reg[165]  ( .D(N9489), .CP(clk), .CD(n3945), .Q(
        mem_data1[165]) );
  CFD2QXL \mem_data1_reg[166]  ( .D(N9490), .CP(clk), .CD(n3946), .Q(
        mem_data1[166]) );
  CFD2QXL \mem_data1_reg[167]  ( .D(N9491), .CP(clk), .CD(n3946), .Q(
        mem_data1[167]) );
  CFD2QXL \mem_data1_reg[168]  ( .D(N9492), .CP(clk), .CD(n3946), .Q(
        mem_data1[168]) );
  CFD2QXL \mem_data1_reg[169]  ( .D(N9493), .CP(clk), .CD(n3946), .Q(
        mem_data1[169]) );
  CFD2QXL \mem_data1_reg[170]  ( .D(N9494), .CP(clk), .CD(n3946), .Q(
        mem_data1[170]) );
  CFD2QXL \mem_data1_reg[171]  ( .D(N9495), .CP(clk), .CD(n3946), .Q(
        mem_data1[171]) );
  CFD2QXL \mem_data1_reg[172]  ( .D(N9496), .CP(clk), .CD(n3946), .Q(
        mem_data1[172]) );
  CFD2QXL \mem_data1_reg[173]  ( .D(N9497), .CP(clk), .CD(n3946), .Q(
        mem_data1[173]) );
  CFD2QXL \mem_data1_reg[174]  ( .D(N9498), .CP(clk), .CD(n3946), .Q(
        mem_data1[174]) );
  CFD2QXL \mem_data1_reg[175]  ( .D(N9499), .CP(clk), .CD(n3946), .Q(
        mem_data1[175]) );
  CFD2QXL \mem_data1_reg[176]  ( .D(N9500), .CP(clk), .CD(n3946), .Q(
        mem_data1[176]) );
  CFD2QXL \mem_data1_reg[177]  ( .D(N9501), .CP(clk), .CD(n3946), .Q(
        mem_data1[177]) );
  CFD2QXL \mem_data1_reg[178]  ( .D(N9502), .CP(clk), .CD(n3946), .Q(
        mem_data1[178]) );
  CFD2QXL \mem_data1_reg[179]  ( .D(N9503), .CP(clk), .CD(n3947), .Q(
        mem_data1[179]) );
  CFD2QXL \mem_data1_reg[180]  ( .D(N9504), .CP(clk), .CD(n3947), .Q(
        mem_data1[180]) );
  CFD2QXL \mem_data1_reg[184]  ( .D(N9508), .CP(clk), .CD(n3947), .Q(
        mem_data1[184]) );
  CFD2QXL \mem_data1_reg[188]  ( .D(N9512), .CP(clk), .CD(n3947), .Q(
        mem_data1[188]) );
  CFD2QXL \mem_data1_reg[190]  ( .D(N9514), .CP(clk), .CD(n3947), .Q(
        mem_data1[190]) );
  CFD2QXL \mem_data1_reg[191]  ( .D(N9515), .CP(clk), .CD(n3947), .Q(
        mem_data1[191]) );
  CFD2QXL \mem_data1_reg[192]  ( .D(N9516), .CP(clk), .CD(n3948), .Q(
        mem_data1[192]) );
  CFD2QXL \mem_data1_reg[193]  ( .D(N9517), .CP(clk), .CD(n3948), .Q(
        mem_data1[193]) );
  CFD2QXL \mem_data1_reg[194]  ( .D(N9518), .CP(clk), .CD(n3948), .Q(
        mem_data1[194]) );
  CFD2QXL \mem_data1_reg[195]  ( .D(N9519), .CP(clk), .CD(n3948), .Q(
        mem_data1[195]) );
  CFD2QXL \mem_data1_reg[196]  ( .D(N9520), .CP(clk), .CD(n3948), .Q(
        mem_data1[196]) );
  CFD2QXL \mem_data1_reg[197]  ( .D(N9521), .CP(clk), .CD(n3948), .Q(
        mem_data1[197]) );
  CFD2QXL \mem_data1_reg[198]  ( .D(N9522), .CP(clk), .CD(n3948), .Q(
        mem_data1[198]) );
  CFD2QXL \mem_data1_reg[199]  ( .D(N9523), .CP(clk), .CD(n3948), .Q(
        mem_data1[199]) );
  CFD2QXL \mem_data1_reg[200]  ( .D(N9524), .CP(clk), .CD(n3948), .Q(
        mem_data1[200]) );
  CFD2QXL \mem_data1_reg[201]  ( .D(N9525), .CP(clk), .CD(n3948), .Q(
        mem_data1[201]) );
  CFD2QXL \mem_data1_reg[202]  ( .D(N9526), .CP(clk), .CD(n3948), .Q(
        mem_data1[202]) );
  CFD2QXL \mem_data1_reg[203]  ( .D(N9527), .CP(clk), .CD(n3948), .Q(
        mem_data1[203]) );
  CFD2QXL \mem_data1_reg[204]  ( .D(N9528), .CP(clk), .CD(n3948), .Q(
        mem_data1[204]) );
  CFD2QXL \mem_data1_reg[205]  ( .D(N9529), .CP(clk), .CD(n3949), .Q(
        mem_data1[205]) );
  CFD2QXL \mem_data1_reg[206]  ( .D(N9530), .CP(clk), .CD(n3949), .Q(
        mem_data1[206]) );
  CFD2QXL \mem_data1_reg[207]  ( .D(N9531), .CP(clk), .CD(n3949), .Q(
        mem_data1[207]) );
  CFD2QXL \mem_data1_reg[208]  ( .D(N9532), .CP(clk), .CD(n3949), .Q(
        mem_data1[208]) );
  CFD2QXL \mem_data1_reg[209]  ( .D(N9533), .CP(clk), .CD(n3949), .Q(
        mem_data1[209]) );
  CFD2QXL \mem_data1_reg[210]  ( .D(N9534), .CP(clk), .CD(n3949), .Q(
        mem_data1[210]) );
  CFD2QXL \mem_data1_reg[211]  ( .D(N9535), .CP(clk), .CD(n3949), .Q(
        mem_data1[211]) );
  CFD2QXL \mem_data1_reg[212]  ( .D(N9536), .CP(clk), .CD(n3949), .Q(
        mem_data1[212]) );
  CFD2QXL \mem_data1_reg[213]  ( .D(N9537), .CP(clk), .CD(n3949), .Q(
        mem_data1[213]) );
  CFD2QXL \mem_data1_reg[214]  ( .D(N9538), .CP(clk), .CD(n3949), .Q(
        mem_data1[214]) );
  CFD2QXL \mem_data1_reg[215]  ( .D(N9539), .CP(clk), .CD(n3949), .Q(
        mem_data1[215]) );
  CFD2QXL \mem_data1_reg[216]  ( .D(N9540), .CP(clk), .CD(n3949), .Q(
        mem_data1[216]) );
  CFD2QXL \mem_data1_reg[217]  ( .D(N9541), .CP(clk), .CD(n3949), .Q(
        mem_data1[217]) );
  CFD2QXL \mem_data1_reg[218]  ( .D(N9542), .CP(clk), .CD(n3950), .Q(
        mem_data1[218]) );
  CFD2QXL \mem_data1_reg[219]  ( .D(N9543), .CP(clk), .CD(n3950), .Q(
        mem_data1[219]) );
  CFD2QXL \mem_data1_reg[221]  ( .D(N9545), .CP(clk), .CD(n3950), .Q(
        mem_data1[221]) );
  CFD2QXL \mem_data1_reg[222]  ( .D(N9546), .CP(clk), .CD(n3950), .Q(
        mem_data1[222]) );
  CFD2QXL \mem_data1_reg[223]  ( .D(N9547), .CP(clk), .CD(n3950), .Q(
        mem_data1[223]) );
  CFD2QXL \mem_data1_reg[224]  ( .D(N9548), .CP(clk), .CD(n3950), .Q(
        mem_data1[224]) );
  CFD2QXL \mem_data1_reg[225]  ( .D(N9549), .CP(clk), .CD(n3976), .Q(
        mem_data1[225]) );
  CFD2QXL \mem_data1_reg[226]  ( .D(N9550), .CP(clk), .CD(n3971), .Q(
        mem_data1[226]) );
  CFD2QXL \mem_data1_reg[229]  ( .D(N9553), .CP(clk), .CD(n3971), .Q(
        mem_data1[229]) );
  CFD2QXL \mem_data1_reg[231]  ( .D(N9555), .CP(clk), .CD(n3971), .Q(
        mem_data1[231]) );
  CFD2QXL \mem_data1_reg[233]  ( .D(N9557), .CP(clk), .CD(n3971), .Q(
        mem_data1[233]) );
  CFD2QXL \mem_data1_reg[235]  ( .D(N9559), .CP(clk), .CD(n3972), .Q(
        mem_data1[235]) );
  CFD2QXL \mem_data1_reg[236]  ( .D(N9560), .CP(clk), .CD(n3972), .Q(
        mem_data1[236]) );
  CFD2QXL \mem_data1_reg[237]  ( .D(N9561), .CP(clk), .CD(n3972), .Q(
        mem_data1[237]) );
  CFD2QXL \mem_data1_reg[240]  ( .D(N9564), .CP(clk), .CD(n3972), .Q(
        mem_data1[240]) );
  CFD2QXL \mem_data1_reg[258]  ( .D(N9582), .CP(clk), .CD(n3973), .Q(
        mem_data1[258]) );
  CFD2QXL \mem_data1_reg[260]  ( .D(N9584), .CP(clk), .CD(n3973), .Q(
        mem_data1[260]) );
  CFD2QXL \mem_data1_reg[262]  ( .D(N9586), .CP(clk), .CD(n3974), .Q(
        mem_data1[262]) );
  CFD2QXL \mem_data1_reg[263]  ( .D(N9587), .CP(clk), .CD(n3974), .Q(
        mem_data1[263]) );
  CFD2QXL \mem_data1_reg[264]  ( .D(N9588), .CP(clk), .CD(n3974), .Q(
        mem_data1[264]) );
  CFD2QXL \mem_data1_reg[265]  ( .D(N9589), .CP(clk), .CD(n3974), .Q(
        mem_data1[265]) );
  CFD2QXL \mem_data1_reg[266]  ( .D(N9590), .CP(clk), .CD(n3974), .Q(
        mem_data1[266]) );
  CFD2QXL \mem_data1_reg[267]  ( .D(N9591), .CP(clk), .CD(n3974), .Q(
        mem_data1[267]) );
  CFD2QXL \mem_data1_reg[268]  ( .D(N9592), .CP(clk), .CD(n3974), .Q(
        mem_data1[268]) );
  CFD2QXL \mem_data1_reg[269]  ( .D(N9593), .CP(clk), .CD(n3974), .Q(
        mem_data1[269]) );
  CFD2QXL \mem_data1_reg[270]  ( .D(N9594), .CP(clk), .CD(n3974), .Q(
        mem_data1[270]) );
  CFD2QXL \mem_data1_reg[272]  ( .D(N9596), .CP(clk), .CD(n3974), .Q(
        mem_data1[272]) );
  CFD2QXL \mem_data1_reg[274]  ( .D(N9598), .CP(clk), .CD(n3975), .Q(
        mem_data1[274]) );
  CFD2QXL \mem_data1_reg[275]  ( .D(N9599), .CP(clk), .CD(n3975), .Q(
        mem_data1[275]) );
  CFD2QXL \mem_data1_reg[276]  ( .D(N9600), .CP(clk), .CD(n3975), .Q(
        mem_data1[276]) );
  CFD2QXL \mem_data1_reg[280]  ( .D(N9604), .CP(clk), .CD(n3975), .Q(
        mem_data1[280]) );
  CFD2QXL \mem_data1_reg[281]  ( .D(N9605), .CP(clk), .CD(n3975), .Q(
        mem_data1[281]) );
  CFD2QXL \mem_data1_reg[284]  ( .D(N9608), .CP(clk), .CD(n3975), .Q(
        mem_data1[284]) );
  CFD2QXL \mem_data1_reg[285]  ( .D(N9609), .CP(clk), .CD(n3975), .Q(
        mem_data1[285]) );
  CFD2QXL \mem_data1_reg[287]  ( .D(N9611), .CP(clk), .CD(n3976), .Q(
        mem_data1[287]) );
  CFD2QXL \mem_data1_reg[288]  ( .D(N9612), .CP(clk), .CD(n3976), .Q(
        mem_data1[288]) );
  CFD2QXL \mem_data1_reg[289]  ( .D(N9613), .CP(clk), .CD(n3976), .Q(
        mem_data1[289]) );
  CFD2QXL \mem_data1_reg[302]  ( .D(N9626), .CP(clk), .CD(n3977), .Q(
        mem_data1[302]) );
  CFD2QXL \mem_data1_reg[306]  ( .D(N9630), .CP(clk), .CD(n3977), .Q(
        mem_data1[306]) );
  CFD2QXL \mem_data1_reg[307]  ( .D(N9631), .CP(clk), .CD(n3977), .Q(
        mem_data1[307]) );
  CFD2QXL \mem_data1_reg[308]  ( .D(N9632), .CP(clk), .CD(n3977), .Q(
        mem_data1[308]) );
  CFD2QXL \mem_data1_reg[310]  ( .D(N9634), .CP(clk), .CD(n3977), .Q(
        mem_data1[310]) );
  CFD2QXL \mem_data1_reg[311]  ( .D(N9635), .CP(clk), .CD(n3977), .Q(
        mem_data1[311]) );
  CFD2QXL \mem_data1_reg[312]  ( .D(N9636), .CP(clk), .CD(n3978), .Q(
        mem_data1[312]) );
  CFD2QXL \mem_data1_reg[318]  ( .D(N9642), .CP(clk), .CD(n3978), .Q(
        mem_data1[318]) );
  CFD2QXL \mem_data1_reg[322]  ( .D(N9646), .CP(clk), .CD(n3978), .Q(
        mem_data1[322]) );
  CFD2QXL \mem_data1_reg[328]  ( .D(N9652), .CP(clk), .CD(n3979), .Q(
        mem_data1[328]) );
  CFD2QXL \mem_data1_reg[329]  ( .D(N9653), .CP(clk), .CD(n3979), .Q(
        mem_data1[329]) );
  CFD2QXL \mem_data1_reg[330]  ( .D(N9654), .CP(clk), .CD(n3979), .Q(
        mem_data1[330]) );
  CFD2QXL \mem_data1_reg[331]  ( .D(N9655), .CP(clk), .CD(n3979), .Q(
        mem_data1[331]) );
  CFD2QXL \mem_data1_reg[332]  ( .D(N9656), .CP(clk), .CD(n3979), .Q(
        mem_data1[332]) );
  CFD2QXL \mem_data1_reg[333]  ( .D(N9657), .CP(clk), .CD(n3979), .Q(
        mem_data1[333]) );
  CFD2QXL \mem_data1_reg[334]  ( .D(N9658), .CP(clk), .CD(n3979), .Q(
        mem_data1[334]) );
  CFD2QXL \mem_data1_reg[336]  ( .D(N9660), .CP(clk), .CD(n3980), .Q(
        mem_data1[336]) );
  CFD2QXL \mem_data1_reg[338]  ( .D(N9662), .CP(clk), .CD(n3980), .Q(
        mem_data1[338]) );
  CFD2QXL \mem_data1_reg[368]  ( .D(N9692), .CP(clk), .CD(n3961), .Q(
        mem_data1[368]) );
  CFD2QXL \mem_data1_reg[382]  ( .D(N9706), .CP(clk), .CD(n3962), .Q(
        mem_data1[382]) );
  CFD2QXL \mem_data1_reg[384]  ( .D(N9708), .CP(clk), .CD(n3962), .Q(
        mem_data1[384]) );
  CFD2QXL \mem_data1_reg[390]  ( .D(N9714), .CP(clk), .CD(n3963), .Q(
        mem_data1[390]) );
  CFD2QXL \mem_data1_reg[392]  ( .D(N9716), .CP(clk), .CD(n3963), .Q(
        mem_data1[392]) );
  CFD2QXL \mem_data1_reg[394]  ( .D(N9718), .CP(clk), .CD(n3963), .Q(
        mem_data1[394]) );
  CFD2QXL \mem_data1_reg[400]  ( .D(N9724), .CP(clk), .CD(n3963), .Q(
        mem_data1[400]) );
  CFD2QXL \mem_data1_reg[403]  ( .D(N9727), .CP(clk), .CD(n3964), .Q(
        mem_data1[403]) );
  CFD2QXL \mem_data1_reg[406]  ( .D(N9730), .CP(clk), .CD(n3964), .Q(
        mem_data1[406]) );
  CFD2QXL \mem_data1_reg[414]  ( .D(N9738), .CP(clk), .CD(n3965), .Q(
        mem_data1[414]) );
  CFD2QXL \mem_data1_reg[420]  ( .D(N9744), .CP(clk), .CD(n3965), .Q(
        mem_data1[420]) );
  CFD2QXL \mem_data1_reg[424]  ( .D(N9748), .CP(clk), .CD(n3965), .Q(
        mem_data1[424]) );
  CFD2QXL \mem_data1_reg[448]  ( .D(N9772), .CP(clk), .CD(n3967), .Q(
        mem_data1[448]) );
  CFD2QXL \mem_data1_reg[449]  ( .D(N9773), .CP(clk), .CD(n3967), .Q(
        mem_data1[449]) );
  CFD2QXL \mem_data1_reg[452]  ( .D(N9776), .CP(clk), .CD(n3968), .Q(
        mem_data1[452]) );
  CFD2QXL \mem_data1_reg[454]  ( .D(N9778), .CP(clk), .CD(n3968), .Q(
        mem_data1[454]) );
  CFD2QXL \mem_data1_reg[456]  ( .D(N9780), .CP(clk), .CD(n3968), .Q(
        mem_data1[456]) );
  CFD2QXL \mem_data1_reg[458]  ( .D(N9782), .CP(clk), .CD(n3968), .Q(
        mem_data1[458]) );
  CFD2QXL \mem_data1_reg[459]  ( .D(N9783), .CP(clk), .CD(n3968), .Q(
        mem_data1[459]) );
  CFD2QXL \mem_data1_reg[462]  ( .D(N9786), .CP(clk), .CD(n3968), .Q(
        mem_data1[462]) );
  CFD2QXL \mem_data1_reg[466]  ( .D(N9790), .CP(clk), .CD(n3969), .Q(
        mem_data1[466]) );
  CFD2QXL \mem_data1_reg[467]  ( .D(N9791), .CP(clk), .CD(n3969), .Q(
        mem_data1[467]) );
  CFD2QXL \mem_data1_reg[468]  ( .D(N9792), .CP(clk), .CD(n3969), .Q(
        mem_data1[468]) );
  CFD2QXL \mem_data1_reg[470]  ( .D(N9794), .CP(clk), .CD(n3969), .Q(
        mem_data1[470]) );
  CFD2QXL \mem_data1_reg[471]  ( .D(N9795), .CP(clk), .CD(n3969), .Q(
        mem_data1[471]) );
  CFD2QXL \mem_data1_reg[472]  ( .D(N9796), .CP(clk), .CD(n3969), .Q(
        mem_data1[472]) );
  CFD2QXL \mem_data1_reg[474]  ( .D(N9798), .CP(clk), .CD(n3969), .Q(
        mem_data1[474]) );
  CFD2QXL \mem_data1_reg[476]  ( .D(N9800), .CP(clk), .CD(n3969), .Q(
        mem_data1[476]) );
  CFD2QXL \mem_data1_reg[478]  ( .D(N9802), .CP(clk), .CD(n3970), .Q(
        mem_data1[478]) );
  CFD2QXL \mem_data1_reg[479]  ( .D(N9803), .CP(clk), .CD(n3970), .Q(
        mem_data1[479]) );
  CFD2QXL \mem_data1_reg[494]  ( .D(N9818), .CP(clk), .CD(n3971), .Q(
        mem_data1[494]) );
  CFD2QXL \mem_data1_reg[497]  ( .D(N9821), .CP(clk), .CD(n3909), .Q(
        mem_data1[497]) );
  CFD2QXL \mem_data1_reg[498]  ( .D(N9822), .CP(clk), .CD(n3909), .Q(
        mem_data1[498]) );
  CFD2QXL \mem_data1_reg[500]  ( .D(N9824), .CP(clk), .CD(n3909), .Q(
        mem_data1[500]) );
  CFD2QXL \mem_data1_reg[501]  ( .D(N9825), .CP(clk), .CD(n3909), .Q(
        mem_data1[501]) );
  CFD2QXL \mem_data1_reg[502]  ( .D(N9826), .CP(clk), .CD(n3909), .Q(
        mem_data1[502]) );
  CFD2QXL \mem_data1_reg[503]  ( .D(N9827), .CP(clk), .CD(n3910), .Q(
        mem_data1[503]) );
  CFD2QXL \mem_data1_reg[504]  ( .D(N9828), .CP(clk), .CD(n3910), .Q(
        mem_data1[504]) );
  CFD2QXL \mem_data1_reg[505]  ( .D(N9829), .CP(clk), .CD(n3910), .Q(
        mem_data1[505]) );
  CFD2QXL \mem_data1_reg[506]  ( .D(N9830), .CP(clk), .CD(n3910), .Q(
        mem_data1[506]) );
  CFD2QXL \mem_data1_reg[507]  ( .D(N9831), .CP(clk), .CD(n3910), .Q(
        mem_data1[507]) );
  CFD2QXL \mem_data1_reg[508]  ( .D(N9832), .CP(clk), .CD(n3910), .Q(
        mem_data1[508]) );
  CFD2QXL \mem_data1_reg[509]  ( .D(N9833), .CP(clk), .CD(n3910), .Q(
        mem_data1[509]) );
  CFD2QXL \mem_data1_reg[510]  ( .D(N9834), .CP(clk), .CD(n3910), .Q(
        mem_data1[510]) );
  CFD2QXL \mem_data1_reg[511]  ( .D(N9835), .CP(clk), .CD(n3910), .Q(
        mem_data1[511]) );
  CFD2QXL \mem_data1_reg[512]  ( .D(N9836), .CP(clk), .CD(n3910), .Q(
        mem_data1[512]) );
  CFD2QXL \mem_data1_reg[513]  ( .D(N9837), .CP(clk), .CD(n3910), .Q(
        mem_data1[513]) );
  CFD2QXL \mem_data1_reg[514]  ( .D(N9838), .CP(clk), .CD(n3910), .Q(
        mem_data1[514]) );
  CFD2QXL \mem_data1_reg[515]  ( .D(N9839), .CP(clk), .CD(n3910), .Q(
        mem_data1[515]) );
  CFD2QXL \mem_data1_reg[516]  ( .D(N9840), .CP(clk), .CD(n3911), .Q(
        mem_data1[516]) );
  CFD2QXL \mem_data1_reg[517]  ( .D(N9841), .CP(clk), .CD(n3911), .Q(
        mem_data1[517]) );
  CFD2QXL \mem_data1_reg[518]  ( .D(N9842), .CP(clk), .CD(n3911), .Q(
        mem_data1[518]) );
  CFD2QXL \mem_data1_reg[519]  ( .D(N9843), .CP(clk), .CD(n3911), .Q(
        mem_data1[519]) );
  CFD2QXL \mem_data1_reg[520]  ( .D(N9844), .CP(clk), .CD(n3911), .Q(
        mem_data1[520]) );
  CFD2QXL \mem_data1_reg[521]  ( .D(N9845), .CP(clk), .CD(n3911), .Q(
        mem_data1[521]) );
  CFD2QXL \mem_data1_reg[522]  ( .D(N9846), .CP(clk), .CD(n3911), .Q(
        mem_data1[522]) );
  CFD2QXL \mem_data1_reg[523]  ( .D(N9847), .CP(clk), .CD(n3911), .Q(
        mem_data1[523]) );
  CFD2QXL \mem_data1_reg[524]  ( .D(N9848), .CP(clk), .CD(n3911), .Q(
        mem_data1[524]) );
  CFD2QXL \mem_data1_reg[525]  ( .D(N9849), .CP(clk), .CD(n3911), .Q(
        mem_data1[525]) );
  CFD2QXL \mem_data1_reg[526]  ( .D(N9850), .CP(clk), .CD(n3911), .Q(
        mem_data1[526]) );
  CFD2QXL \mem_data1_reg[527]  ( .D(N9851), .CP(clk), .CD(n3911), .Q(
        mem_data1[527]) );
  CFD2QXL \mem_data1_reg[528]  ( .D(N9852), .CP(clk), .CD(n3911), .Q(
        mem_data1[528]) );
  CFD2QXL \mem_data1_reg[529]  ( .D(N9853), .CP(clk), .CD(n3912), .Q(
        mem_data1[529]) );
  CFD2QXL \mem_data1_reg[530]  ( .D(N9854), .CP(clk), .CD(n3912), .Q(
        mem_data1[530]) );
  CFD2QXL \mem_data1_reg[531]  ( .D(N9855), .CP(clk), .CD(n3912), .Q(
        mem_data1[531]) );
  CFD2QXL \mem_data1_reg[532]  ( .D(N9856), .CP(clk), .CD(n3912), .Q(
        mem_data1[532]) );
  CFD2QXL \mem_data1_reg[533]  ( .D(N9857), .CP(clk), .CD(n3912), .Q(
        mem_data1[533]) );
  CFD2QXL \mem_data1_reg[534]  ( .D(N9858), .CP(clk), .CD(n3912), .Q(
        mem_data1[534]) );
  CFD2QXL \mem_data1_reg[535]  ( .D(N9859), .CP(clk), .CD(n3912), .Q(
        mem_data1[535]) );
  CFD2QXL \mem_data1_reg[536]  ( .D(N9860), .CP(clk), .CD(n3912), .Q(
        mem_data1[536]) );
  CFD2QXL \mem_data1_reg[537]  ( .D(N9861), .CP(clk), .CD(n3912), .Q(
        mem_data1[537]) );
  CFD2QXL \mem_data1_reg[538]  ( .D(N9862), .CP(clk), .CD(n3912), .Q(
        mem_data1[538]) );
  CFD2QXL \mem_data1_reg[539]  ( .D(N9863), .CP(clk), .CD(n3912), .Q(
        mem_data1[539]) );
  CFD2QXL \mem_data1_reg[540]  ( .D(N9864), .CP(clk), .CD(n3912), .Q(
        mem_data1[540]) );
  CFD2QXL \mem_data1_reg[541]  ( .D(N9865), .CP(clk), .CD(n3912), .Q(
        mem_data1[541]) );
  CFD2QXL \mem_data1_reg[542]  ( .D(N9866), .CP(clk), .CD(n3913), .Q(
        mem_data1[542]) );
  CFD2QXL \mem_data1_reg[543]  ( .D(N9867), .CP(clk), .CD(n3913), .Q(
        mem_data1[543]) );
  CFD2QXL \mem_data1_reg[544]  ( .D(N9868), .CP(clk), .CD(n3913), .Q(
        mem_data1[544]) );
  CFD2QXL \mem_data1_reg[545]  ( .D(N9869), .CP(clk), .CD(n3913), .Q(
        mem_data1[545]) );
  CFD2QXL \mem_data1_reg[546]  ( .D(N9870), .CP(clk), .CD(n3913), .Q(
        mem_data1[546]) );
  CFD2QXL \mem_data1_reg[547]  ( .D(N9871), .CP(clk), .CD(n3913), .Q(
        mem_data1[547]) );
  CFD2QXL \mem_data1_reg[548]  ( .D(N9872), .CP(clk), .CD(n3913), .Q(
        mem_data1[548]) );
  CFD2QXL \mem_data1_reg[549]  ( .D(N9873), .CP(clk), .CD(n3913), .Q(
        mem_data1[549]) );
  CFD2QXL \mem_data1_reg[550]  ( .D(N9874), .CP(clk), .CD(n3913), .Q(
        mem_data1[550]) );
  CFD2QXL \mem_data1_reg[551]  ( .D(N9875), .CP(clk), .CD(n3913), .Q(
        mem_data1[551]) );
  CFD2QXL \mem_data1_reg[552]  ( .D(N9876), .CP(clk), .CD(n3913), .Q(
        mem_data1[552]) );
  CFD2QXL \mem_data1_reg[553]  ( .D(N9877), .CP(clk), .CD(n3913), .Q(
        mem_data1[553]) );
  CFD2QXL \mem_data1_reg[554]  ( .D(N9878), .CP(clk), .CD(n3913), .Q(
        mem_data1[554]) );
  CFD2QXL \mem_data1_reg[555]  ( .D(N9879), .CP(clk), .CD(n3914), .Q(
        mem_data1[555]) );
  CFD2QXL \mem_data1_reg[556]  ( .D(N9880), .CP(clk), .CD(n3914), .Q(
        mem_data1[556]) );
  CFD2QXL \mem_data1_reg[557]  ( .D(N9881), .CP(clk), .CD(n3914), .Q(
        mem_data1[557]) );
  CFD2QXL \mem_data1_reg[558]  ( .D(N9882), .CP(clk), .CD(n3914), .Q(
        mem_data1[558]) );
  CFD2QXL \mem_data1_reg[559]  ( .D(N9883), .CP(clk), .CD(n3914), .Q(
        mem_data1[559]) );
  CFD2QXL \mem_data1_reg[560]  ( .D(N9884), .CP(clk), .CD(n3914), .Q(
        mem_data1[560]) );
  CFD2QXL \mem_data1_reg[561]  ( .D(N9885), .CP(clk), .CD(n3914), .Q(
        mem_data1[561]) );
  CFD2QXL \mem_data1_reg[562]  ( .D(N9886), .CP(clk), .CD(n3914), .Q(
        mem_data1[562]) );
  CFD2QXL \mem_data1_reg[563]  ( .D(N9887), .CP(clk), .CD(n3914), .Q(
        mem_data1[563]) );
  CFD2QXL \mem_data1_reg[564]  ( .D(N9888), .CP(clk), .CD(n3914), .Q(
        mem_data1[564]) );
  CFD2QXL \mem_data1_reg[565]  ( .D(N9889), .CP(clk), .CD(n3914), .Q(
        mem_data1[565]) );
  CFD2QXL \mem_data1_reg[566]  ( .D(N9890), .CP(clk), .CD(n3914), .Q(
        mem_data1[566]) );
  CFD2QXL \mem_data1_reg[567]  ( .D(N9891), .CP(clk), .CD(n3915), .Q(
        mem_data1[567]) );
  CFD2QXL \mem_data1_reg[568]  ( .D(N9892), .CP(clk), .CD(n3915), .Q(
        mem_data1[568]) );
  CFD2QXL \mem_data1_reg[569]  ( .D(N9893), .CP(clk), .CD(n3915), .Q(
        mem_data1[569]) );
  CFD2QXL \mem_data1_reg[570]  ( .D(N9894), .CP(clk), .CD(n3915), .Q(
        mem_data1[570]) );
  CFD2QXL \mem_data1_reg[571]  ( .D(N9895), .CP(clk), .CD(n3915), .Q(
        mem_data1[571]) );
  CFD2QXL \mem_data1_reg[572]  ( .D(N9896), .CP(clk), .CD(n3915), .Q(
        mem_data1[572]) );
  CFD2QXL \mem_data1_reg[573]  ( .D(N9897), .CP(clk), .CD(n3915), .Q(
        mem_data1[573]) );
  CFD2QXL \mem_data1_reg[574]  ( .D(N9898), .CP(clk), .CD(n3915), .Q(
        mem_data1[574]) );
  CFD2QXL \mem_data1_reg[575]  ( .D(N9899), .CP(clk), .CD(n3915), .Q(
        mem_data1[575]) );
  CFD2QXL \mem_data1_reg[576]  ( .D(N9900), .CP(clk), .CD(n3915), .Q(
        mem_data1[576]) );
  CFD2QXL \mem_data1_reg[577]  ( .D(N9901), .CP(clk), .CD(n3915), .Q(
        mem_data1[577]) );
  CFD2QXL \mem_data1_reg[578]  ( .D(N9902), .CP(clk), .CD(n3915), .Q(
        mem_data1[578]) );
  CFD2QXL \mem_data1_reg[579]  ( .D(N9903), .CP(clk), .CD(n3915), .Q(
        mem_data1[579]) );
  CFD2QXL \mem_data1_reg[580]  ( .D(N9904), .CP(clk), .CD(n3916), .Q(
        mem_data1[580]) );
  CFD2QXL \mem_data1_reg[581]  ( .D(N9905), .CP(clk), .CD(n3916), .Q(
        mem_data1[581]) );
  CFD2QXL \mem_data1_reg[582]  ( .D(N9906), .CP(clk), .CD(n3916), .Q(
        mem_data1[582]) );
  CFD2QXL \mem_data1_reg[583]  ( .D(N9907), .CP(clk), .CD(n3916), .Q(
        mem_data1[583]) );
  CFD2QXL \mem_data1_reg[584]  ( .D(N9908), .CP(clk), .CD(n3916), .Q(
        mem_data1[584]) );
  CFD2QXL \mem_data1_reg[585]  ( .D(N9909), .CP(clk), .CD(n3916), .Q(
        mem_data1[585]) );
  CFD2QXL \mem_data1_reg[586]  ( .D(N9910), .CP(clk), .CD(n3916), .Q(
        mem_data1[586]) );
  CFD2QXL \mem_data1_reg[587]  ( .D(N9911), .CP(clk), .CD(n3916), .Q(
        mem_data1[587]) );
  CFD2QXL \mem_data1_reg[588]  ( .D(N9912), .CP(clk), .CD(n3916), .Q(
        mem_data1[588]) );
  CFD2QXL \mem_data1_reg[589]  ( .D(N9913), .CP(clk), .CD(n3916), .Q(
        mem_data1[589]) );
  CFD2QXL \mem_data1_reg[590]  ( .D(N9914), .CP(clk), .CD(n3916), .Q(
        mem_data1[590]) );
  CFD2QXL \mem_data1_reg[591]  ( .D(N9915), .CP(clk), .CD(n3916), .Q(
        mem_data1[591]) );
  CFD2QXL \mem_data1_reg[592]  ( .D(N9916), .CP(clk), .CD(n3916), .Q(
        mem_data1[592]) );
  CFD2QXL \mem_data1_reg[593]  ( .D(N9917), .CP(clk), .CD(n3917), .Q(
        mem_data1[593]) );
  CFD2QXL \mem_data1_reg[594]  ( .D(N9918), .CP(clk), .CD(n3917), .Q(
        mem_data1[594]) );
  CFD2QXL \mem_data1_reg[595]  ( .D(N9919), .CP(clk), .CD(n3917), .Q(
        mem_data1[595]) );
  CFD2QXL \mem_data1_reg[596]  ( .D(N9920), .CP(clk), .CD(n3917), .Q(
        mem_data1[596]) );
  CFD2QXL \mem_data1_reg[597]  ( .D(N9921), .CP(clk), .CD(n3917), .Q(
        mem_data1[597]) );
  CFD2QXL \mem_data1_reg[598]  ( .D(N9922), .CP(clk), .CD(n3917), .Q(
        mem_data1[598]) );
  CFD2QXL \mem_data1_reg[599]  ( .D(N9923), .CP(clk), .CD(n3917), .Q(
        mem_data1[599]) );
  CFD2QXL \mem_data1_reg[600]  ( .D(N9924), .CP(clk), .CD(n3917), .Q(
        mem_data1[600]) );
  CFD2QXL \mem_data1_reg[601]  ( .D(N9925), .CP(clk), .CD(n3917), .Q(
        mem_data1[601]) );
  CFD2QXL \mem_data1_reg[602]  ( .D(N9926), .CP(clk), .CD(n3917), .Q(
        mem_data1[602]) );
  CFD2QXL \mem_data1_reg[603]  ( .D(N9927), .CP(clk), .CD(n3917), .Q(
        mem_data1[603]) );
  CFD2QXL \mem_data1_reg[604]  ( .D(N9928), .CP(clk), .CD(n3917), .Q(
        mem_data1[604]) );
  CFD2QXL \mem_data1_reg[605]  ( .D(N9929), .CP(clk), .CD(n3917), .Q(
        mem_data1[605]) );
  CFD2QXL \mem_data1_reg[606]  ( .D(N9930), .CP(clk), .CD(n3918), .Q(
        mem_data1[606]) );
  CFD2QXL \mem_data1_reg[607]  ( .D(N9931), .CP(clk), .CD(n3918), .Q(
        mem_data1[607]) );
  CFD2QXL \mem_data1_reg[608]  ( .D(N9932), .CP(clk), .CD(n3918), .Q(
        mem_data1[608]) );
  CFD2QXL \mem_data1_reg[609]  ( .D(N9933), .CP(clk), .CD(n3918), .Q(
        mem_data1[609]) );
  CFD2QXL \mem_data1_reg[610]  ( .D(N9934), .CP(clk), .CD(n3918), .Q(
        mem_data1[610]) );
  CFD2QXL \mem_data1_reg[611]  ( .D(N9935), .CP(clk), .CD(n3918), .Q(
        mem_data1[611]) );
  CFD2QXL \mem_data1_reg[612]  ( .D(N9936), .CP(clk), .CD(n3918), .Q(
        mem_data1[612]) );
  CFD2QXL \mem_data1_reg[613]  ( .D(N9937), .CP(clk), .CD(n3918), .Q(
        mem_data1[613]) );
  CFD2QXL \mem_data1_reg[614]  ( .D(N9938), .CP(clk), .CD(n3918), .Q(
        mem_data1[614]) );
  CFD2QXL \mem_data1_reg[615]  ( .D(N9939), .CP(clk), .CD(n3918), .Q(
        mem_data1[615]) );
  CFD2QXL \mem_data1_reg[616]  ( .D(N9940), .CP(clk), .CD(n3918), .Q(
        mem_data1[616]) );
  CFD2QXL \mem_data1_reg[617]  ( .D(N9941), .CP(clk), .CD(n3918), .Q(
        mem_data1[617]) );
  CFD2QXL \mem_data1_reg[618]  ( .D(N9942), .CP(clk), .CD(n3918), .Q(
        mem_data1[618]) );
  CFD2QXL \mem_data1_reg[619]  ( .D(N9943), .CP(clk), .CD(n3919), .Q(
        mem_data1[619]) );
  CFD2QXL \mem_data1_reg[620]  ( .D(N9944), .CP(clk), .CD(n3919), .Q(
        mem_data1[620]) );
  CFD2QXL \mem_data1_reg[621]  ( .D(N9945), .CP(clk), .CD(n3919), .Q(
        mem_data1[621]) );
  CFD2QXL \mem_data1_reg[622]  ( .D(N9946), .CP(clk), .CD(n3919), .Q(
        mem_data1[622]) );
  CFD2QXL \mem_data1_reg[623]  ( .D(N9947), .CP(clk), .CD(n3919), .Q(
        mem_data1[623]) );
  CFD2QXL \mem_data1_reg[624]  ( .D(N9948), .CP(clk), .CD(n3919), .Q(
        mem_data1[624]) );
  CFD2QXL \mem_data1_reg[625]  ( .D(N9949), .CP(clk), .CD(n3919), .Q(
        mem_data1[625]) );
  CFD2QXL \mem_data1_reg[626]  ( .D(N9950), .CP(clk), .CD(n3919), .Q(
        mem_data1[626]) );
  CFD2QXL \mem_data1_reg[627]  ( .D(N9951), .CP(clk), .CD(n3919), .Q(
        mem_data1[627]) );
  CFD2QXL \mem_data1_reg[628]  ( .D(N9952), .CP(clk), .CD(n3904), .Q(
        mem_data1[628]) );
  CFD2QXL \mem_data1_reg[629]  ( .D(N9953), .CP(clk), .CD(n3899), .Q(
        mem_data1[629]) );
  CFD2QXL \mem_data1_reg[630]  ( .D(N9954), .CP(clk), .CD(n3899), .Q(
        mem_data1[630]) );
  CFD2QXL \mem_data1_reg[631]  ( .D(N9955), .CP(clk), .CD(n3899), .Q(
        mem_data1[631]) );
  CFD2QXL \mem_data1_reg[632]  ( .D(N9956), .CP(clk), .CD(n3899), .Q(
        mem_data1[632]) );
  CFD2QXL \mem_data1_reg[633]  ( .D(N9957), .CP(clk), .CD(n3899), .Q(
        mem_data1[633]) );
  CFD2QXL \mem_data1_reg[634]  ( .D(N9958), .CP(clk), .CD(n3899), .Q(
        mem_data1[634]) );
  CFD2QXL \mem_data1_reg[635]  ( .D(N9959), .CP(clk), .CD(n3899), .Q(
        mem_data1[635]) );
  CFD2QXL \mem_data1_reg[636]  ( .D(N9960), .CP(clk), .CD(n3899), .Q(
        mem_data1[636]) );
  CFD2QXL \mem_data1_reg[637]  ( .D(N9961), .CP(clk), .CD(n3900), .Q(
        mem_data1[637]) );
  CFD2QXL \mem_data1_reg[638]  ( .D(N9962), .CP(clk), .CD(n3900), .Q(
        mem_data1[638]) );
  CFD2QXL \mem_data1_reg[639]  ( .D(N9963), .CP(clk), .CD(n3900), .Q(
        mem_data1[639]) );
  CFD2QXL \mem_data1_reg[640]  ( .D(N9964), .CP(clk), .CD(n3900), .Q(
        mem_data1[640]) );
  CFD2QXL \mem_data1_reg[641]  ( .D(N9965), .CP(clk), .CD(n3900), .Q(
        mem_data1[641]) );
  CFD2QXL \mem_data1_reg[642]  ( .D(N9966), .CP(clk), .CD(n3900), .Q(
        mem_data1[642]) );
  CFD2QXL \mem_data1_reg[643]  ( .D(N9967), .CP(clk), .CD(n3900), .Q(
        mem_data1[643]) );
  CFD2QXL \mem_data1_reg[644]  ( .D(N9968), .CP(clk), .CD(n3900), .Q(
        mem_data1[644]) );
  CFD2QXL \mem_data1_reg[645]  ( .D(N9969), .CP(clk), .CD(n3900), .Q(
        mem_data1[645]) );
  CFD2QXL \mem_data1_reg[646]  ( .D(N9970), .CP(clk), .CD(n3900), .Q(
        mem_data1[646]) );
  CFD2QXL \mem_data1_reg[647]  ( .D(N9971), .CP(clk), .CD(n3900), .Q(
        mem_data1[647]) );
  CFD2QXL \mem_data1_reg[648]  ( .D(N9972), .CP(clk), .CD(n3900), .Q(
        mem_data1[648]) );
  CFD2QXL \mem_data1_reg[649]  ( .D(N9973), .CP(clk), .CD(n3900), .Q(
        mem_data1[649]) );
  CFD2QXL \mem_data1_reg[650]  ( .D(N9974), .CP(clk), .CD(n3901), .Q(
        mem_data1[650]) );
  CFD2QXL \mem_data1_reg[651]  ( .D(N9975), .CP(clk), .CD(n3901), .Q(
        mem_data1[651]) );
  CFD2QXL \mem_data1_reg[652]  ( .D(N9976), .CP(clk), .CD(n3901), .Q(
        mem_data1[652]) );
  CFD2QXL \mem_data1_reg[653]  ( .D(N9977), .CP(clk), .CD(n3901), .Q(
        mem_data1[653]) );
  CFD2QXL \mem_data1_reg[654]  ( .D(N9978), .CP(clk), .CD(n3901), .Q(
        mem_data1[654]) );
  CFD2QXL \mem_data1_reg[655]  ( .D(N9979), .CP(clk), .CD(n3901), .Q(
        mem_data1[655]) );
  CFD2QXL \mem_data1_reg[656]  ( .D(N9980), .CP(clk), .CD(n3901), .Q(
        mem_data1[656]) );
  CFD2QXL \mem_data1_reg[657]  ( .D(N9981), .CP(clk), .CD(n3901), .Q(
        mem_data1[657]) );
  CFD2QXL \mem_data1_reg[658]  ( .D(N9982), .CP(clk), .CD(n3901), .Q(
        mem_data1[658]) );
  CFD2QXL \mem_data1_reg[659]  ( .D(N9983), .CP(clk), .CD(n3901), .Q(
        mem_data1[659]) );
  CFD2QXL \mem_data1_reg[660]  ( .D(N9984), .CP(clk), .CD(n3901), .Q(
        mem_data1[660]) );
  CFD2QXL \mem_data1_reg[661]  ( .D(N9985), .CP(clk), .CD(n3901), .Q(
        mem_data1[661]) );
  CFD2QXL \mem_data1_reg[662]  ( .D(N9986), .CP(clk), .CD(n3901), .Q(
        mem_data1[662]) );
  CFD2QXL \mem_data1_reg[663]  ( .D(N9987), .CP(clk), .CD(n3902), .Q(
        mem_data1[663]) );
  CFD2QXL \mem_data1_reg[664]  ( .D(N9988), .CP(clk), .CD(n3902), .Q(
        mem_data1[664]) );
  CFD2QXL \mem_data1_reg[665]  ( .D(N9989), .CP(clk), .CD(n3902), .Q(
        mem_data1[665]) );
  CFD2QXL \mem_data1_reg[666]  ( .D(N9990), .CP(clk), .CD(n3902), .Q(
        mem_data1[666]) );
  CFD2QXL \mem_data1_reg[667]  ( .D(N9991), .CP(clk), .CD(n3902), .Q(
        mem_data1[667]) );
  CFD2QXL \mem_data1_reg[668]  ( .D(N9992), .CP(clk), .CD(n3902), .Q(
        mem_data1[668]) );
  CFD2QXL \mem_data1_reg[669]  ( .D(N9993), .CP(clk), .CD(n3902), .Q(
        mem_data1[669]) );
  CFD2QXL \mem_data1_reg[670]  ( .D(N9994), .CP(clk), .CD(n3902), .Q(
        mem_data1[670]) );
  CFD2QXL \mem_data1_reg[671]  ( .D(N9995), .CP(clk), .CD(n3902), .Q(
        mem_data1[671]) );
  CFD2QXL \mem_data1_reg[672]  ( .D(N9996), .CP(clk), .CD(n3902), .Q(
        mem_data1[672]) );
  CFD2QXL \mem_data1_reg[673]  ( .D(N9997), .CP(clk), .CD(n3902), .Q(
        mem_data1[673]) );
  CFD2QXL \mem_data1_reg[674]  ( .D(N9998), .CP(clk), .CD(n3902), .Q(
        mem_data1[674]) );
  CFD2QXL \mem_data1_reg[675]  ( .D(N9999), .CP(clk), .CD(n3902), .Q(
        mem_data1[675]) );
  CFD2QXL \mem_data1_reg[677]  ( .D(N10001), .CP(clk), .CD(n3903), .Q(
        mem_data1[677]) );
  CFD2QXL \mem_data1_reg[678]  ( .D(N10002), .CP(clk), .CD(n3903), .Q(
        mem_data1[678]) );
  CFD2QXL \mem_data1_reg[679]  ( .D(N10003), .CP(clk), .CD(n3903), .Q(
        mem_data1[679]) );
  CFD2QXL \mem_data1_reg[680]  ( .D(N10004), .CP(clk), .CD(n3903), .Q(
        mem_data1[680]) );
  CFD2QXL \mem_data1_reg[681]  ( .D(N10005), .CP(clk), .CD(n3903), .Q(
        mem_data1[681]) );
  CFD2QXL \mem_data1_reg[682]  ( .D(N10006), .CP(clk), .CD(n3903), .Q(
        mem_data1[682]) );
  CFD2QXL \mem_data1_reg[683]  ( .D(N10007), .CP(clk), .CD(n3903), .Q(
        mem_data1[683]) );
  CFD2QXL \mem_data1_reg[684]  ( .D(N10008), .CP(clk), .CD(n3903), .Q(
        mem_data1[684]) );
  CFD2QXL \mem_data1_reg[685]  ( .D(N10009), .CP(clk), .CD(n3903), .Q(
        mem_data1[685]) );
  CFD2QXL \mem_data1_reg[686]  ( .D(N10010), .CP(clk), .CD(n3903), .Q(
        mem_data1[686]) );
  CFD2QXL \mem_data1_reg[687]  ( .D(N10011), .CP(clk), .CD(n3903), .Q(
        mem_data1[687]) );
  CFD2QXL \mem_data1_reg[688]  ( .D(N10012), .CP(clk), .CD(n3903), .Q(
        mem_data1[688]) );
  CFD2QXL \mem_data1_reg[689]  ( .D(N10013), .CP(clk), .CD(n3903), .Q(
        mem_data1[689]) );
  CFD2QXL \mem_data1_reg[690]  ( .D(N10014), .CP(clk), .CD(n3904), .Q(
        mem_data1[690]) );
  CFD2QXL \mem_data1_reg[691]  ( .D(N10015), .CP(clk), .CD(n3904), .Q(
        mem_data1[691]) );
  CFD2QXL \mem_data1_reg[692]  ( .D(N10016), .CP(clk), .CD(n3904), .Q(
        mem_data1[692]) );
  CFD2QXL \mem_data1_reg[693]  ( .D(N10017), .CP(clk), .CD(n3904), .Q(
        mem_data1[693]) );
  CFD2QXL \mem_data1_reg[694]  ( .D(N10018), .CP(clk), .CD(n3904), .Q(
        mem_data1[694]) );
  CFD2QXL \mem_data1_reg[695]  ( .D(N10019), .CP(clk), .CD(n3904), .Q(
        mem_data1[695]) );
  CFD2QXL \mem_data1_reg[696]  ( .D(N10020), .CP(clk), .CD(n3904), .Q(
        mem_data1[696]) );
  CFD2QXL \mem_data1_reg[697]  ( .D(N10021), .CP(clk), .CD(n3904), .Q(
        mem_data1[697]) );
  CFD2QXL \mem_data1_reg[698]  ( .D(N10022), .CP(clk), .CD(n3904), .Q(
        mem_data1[698]) );
  CFD2QXL \mem_data1_reg[699]  ( .D(N10023), .CP(clk), .CD(n3904), .Q(
        mem_data1[699]) );
  CFD2QXL \mem_data1_reg[700]  ( .D(N10024), .CP(clk), .CD(n3904), .Q(
        mem_data1[700]) );
  CFD2QXL \mem_data1_reg[701]  ( .D(N10025), .CP(clk), .CD(n3904), .Q(
        mem_data1[701]) );
  CFD2QXL \mem_data1_reg[702]  ( .D(N10026), .CP(clk), .CD(n3905), .Q(
        mem_data1[702]) );
  CFD2QXL \mem_data1_reg[703]  ( .D(N10027), .CP(clk), .CD(n3905), .Q(
        mem_data1[703]) );
  CFD2QXL \mem_data1_reg[704]  ( .D(N10028), .CP(clk), .CD(n3905), .Q(
        mem_data1[704]) );
  CFD2QXL \mem_data1_reg[705]  ( .D(N10029), .CP(clk), .CD(n3905), .Q(
        mem_data1[705]) );
  CFD2QXL \mem_data1_reg[706]  ( .D(N10030), .CP(clk), .CD(n3905), .Q(
        mem_data1[706]) );
  CFD2QXL \mem_data1_reg[707]  ( .D(N10031), .CP(clk), .CD(n3905), .Q(
        mem_data1[707]) );
  CFD2QXL \mem_data1_reg[708]  ( .D(N10032), .CP(clk), .CD(n3905), .Q(
        mem_data1[708]) );
  CFD2QXL \mem_data1_reg[709]  ( .D(N10033), .CP(clk), .CD(n3905), .Q(
        mem_data1[709]) );
  CFD2QXL \mem_data1_reg[710]  ( .D(N10034), .CP(clk), .CD(n3905), .Q(
        mem_data1[710]) );
  CFD2QXL \mem_data1_reg[711]  ( .D(N10035), .CP(clk), .CD(n3905), .Q(
        mem_data1[711]) );
  CFD2QXL \mem_data1_reg[712]  ( .D(N10036), .CP(clk), .CD(n3905), .Q(
        mem_data1[712]) );
  CFD2QXL \mem_data1_reg[713]  ( .D(N10037), .CP(clk), .CD(n3905), .Q(
        mem_data1[713]) );
  CFD2QXL \mem_data1_reg[714]  ( .D(N10038), .CP(clk), .CD(n3905), .Q(
        mem_data1[714]) );
  CFD2QXL \mem_data1_reg[715]  ( .D(N10039), .CP(clk), .CD(n3906), .Q(
        mem_data1[715]) );
  CFD2QXL \mem_data1_reg[716]  ( .D(N10040), .CP(clk), .CD(n3906), .Q(
        mem_data1[716]) );
  CFD2QXL \mem_data1_reg[717]  ( .D(N10041), .CP(clk), .CD(n3906), .Q(
        mem_data1[717]) );
  CFD2QXL \mem_data1_reg[718]  ( .D(N10042), .CP(clk), .CD(n3906), .Q(
        mem_data1[718]) );
  CFD2QXL \mem_data1_reg[719]  ( .D(N10043), .CP(clk), .CD(n3906), .Q(
        mem_data1[719]) );
  CFD2QXL \mem_data1_reg[720]  ( .D(N10044), .CP(clk), .CD(n3906), .Q(
        mem_data1[720]) );
  CFD2QXL \mem_data1_reg[721]  ( .D(N10045), .CP(clk), .CD(n3906), .Q(
        mem_data1[721]) );
  CFD2QXL \mem_data1_reg[722]  ( .D(N10046), .CP(clk), .CD(n3906), .Q(
        mem_data1[722]) );
  CFD2QXL \mem_data1_reg[723]  ( .D(N10047), .CP(clk), .CD(n3906), .Q(
        mem_data1[723]) );
  CFD2QXL \mem_data1_reg[724]  ( .D(N10048), .CP(clk), .CD(n3906), .Q(
        mem_data1[724]) );
  CFD2QXL \mem_data1_reg[725]  ( .D(N10049), .CP(clk), .CD(n3906), .Q(
        mem_data1[725]) );
  CFD2QXL \mem_data1_reg[726]  ( .D(N10050), .CP(clk), .CD(n3906), .Q(
        mem_data1[726]) );
  CFD2QXL \mem_data1_reg[727]  ( .D(N10051), .CP(clk), .CD(n3906), .Q(
        mem_data1[727]) );
  CFD2QXL \mem_data1_reg[728]  ( .D(N10052), .CP(clk), .CD(n3907), .Q(
        mem_data1[728]) );
  CFD2QXL \mem_data1_reg[729]  ( .D(N10053), .CP(clk), .CD(n3907), .Q(
        mem_data1[729]) );
  CFD2QXL \mem_data1_reg[730]  ( .D(N10054), .CP(clk), .CD(n3907), .Q(
        mem_data1[730]) );
  CFD2QXL \mem_data1_reg[731]  ( .D(N10055), .CP(clk), .CD(n3907), .Q(
        mem_data1[731]) );
  CFD2QXL \mem_data1_reg[732]  ( .D(N10056), .CP(clk), .CD(n3907), .Q(
        mem_data1[732]) );
  CFD2QXL \mem_data1_reg[733]  ( .D(N10057), .CP(clk), .CD(n3907), .Q(
        mem_data1[733]) );
  CFD2QXL \mem_data1_reg[734]  ( .D(N10058), .CP(clk), .CD(n3907), .Q(
        mem_data1[734]) );
  CFD2QXL \mem_data1_reg[735]  ( .D(N10059), .CP(clk), .CD(n3907), .Q(
        mem_data1[735]) );
  CFD2QXL \mem_data1_reg[736]  ( .D(N10060), .CP(clk), .CD(n3907), .Q(
        mem_data1[736]) );
  CFD2QXL \mem_data1_reg[737]  ( .D(N10061), .CP(clk), .CD(n3907), .Q(
        mem_data1[737]) );
  CFD2QXL \mem_data1_reg[738]  ( .D(N10062), .CP(clk), .CD(n3907), .Q(
        mem_data1[738]) );
  CFD2QXL \mem_data1_reg[739]  ( .D(N10063), .CP(clk), .CD(n3907), .Q(
        mem_data1[739]) );
  CFD2QXL \mem_data1_reg[740]  ( .D(N10064), .CP(clk), .CD(n3907), .Q(
        mem_data1[740]) );
  CFD2QXL \mem_data1_reg[741]  ( .D(N10065), .CP(clk), .CD(n3908), .Q(
        mem_data1[741]) );
  CFD2QXL \mem_data1_reg[742]  ( .D(N10066), .CP(clk), .CD(n3908), .Q(
        mem_data1[742]) );
  CFD2QXL \mem_data1_reg[743]  ( .D(N10067), .CP(clk), .CD(n3908), .Q(
        mem_data1[743]) );
  CFD2QXL \mem_data1_reg[744]  ( .D(N10068), .CP(clk), .CD(n3908), .Q(
        mem_data1[744]) );
  CFD2QXL \mem_data1_reg[745]  ( .D(N10069), .CP(clk), .CD(n3908), .Q(
        mem_data1[745]) );
  CFD2QXL \mem_data1_reg[746]  ( .D(N10070), .CP(clk), .CD(n3908), .Q(
        mem_data1[746]) );
  CFD2QXL \mem_data1_reg[747]  ( .D(N10071), .CP(clk), .CD(n3908), .Q(
        mem_data1[747]) );
  CFD2QXL \mem_data1_reg[748]  ( .D(N10072), .CP(clk), .CD(n3908), .Q(
        mem_data1[748]) );
  CFD2QXL \mem_data1_reg[749]  ( .D(N10073), .CP(clk), .CD(n3908), .Q(
        mem_data1[749]) );
  CFD2QXL \mem_data1_reg[750]  ( .D(N10074), .CP(clk), .CD(n3908), .Q(
        mem_data1[750]) );
  CFD2QXL \mem_data1_reg[751]  ( .D(N10075), .CP(clk), .CD(n3908), .Q(
        mem_data1[751]) );
  CFD2QXL \mem_data1_reg[752]  ( .D(N10076), .CP(clk), .CD(n3908), .Q(
        mem_data1[752]) );
  CFD2QXL \mem_data1_reg[753]  ( .D(N10077), .CP(clk), .CD(n3908), .Q(
        mem_data1[753]) );
  CFD2QXL \mem_data1_reg[754]  ( .D(N10078), .CP(clk), .CD(n3909), .Q(
        mem_data1[754]) );
  CFD2QXL \mem_data1_reg[755]  ( .D(N10079), .CP(clk), .CD(n3909), .Q(
        mem_data1[755]) );
  CFD2QXL \mem_data1_reg[756]  ( .D(N10080), .CP(clk), .CD(n3909), .Q(
        mem_data1[756]) );
  CFD2QXL \mem_data1_reg[757]  ( .D(N10081), .CP(clk), .CD(n3909), .Q(
        mem_data1[757]) );
  CFD2QXL \mem_data1_reg[758]  ( .D(N10082), .CP(clk), .CD(n3909), .Q(
        mem_data1[758]) );
  CFD2QXL \mem_data1_reg[759]  ( .D(N10083), .CP(clk), .CD(n3909), .Q(
        mem_data1[759]) );
  CFD2QXL \mem_data1_reg[760]  ( .D(N10084), .CP(clk), .CD(n3909), .Q(
        mem_data1[760]) );
  CFD2QXL \mem_data1_reg[761]  ( .D(N10085), .CP(clk), .CD(n3934), .Q(
        mem_data1[761]) );
  CFD2QXL \mem_data1_reg[762]  ( .D(N10086), .CP(clk), .CD(n3929), .Q(
        mem_data1[762]) );
  CFD2QXL \mem_data1_reg[763]  ( .D(N10087), .CP(clk), .CD(n3930), .Q(
        mem_data1[763]) );
  CFD2QXL \mem_data1_reg[764]  ( .D(N10088), .CP(clk), .CD(n3930), .Q(
        mem_data1[764]) );
  CFD2QXL \mem_data1_reg[765]  ( .D(N10089), .CP(clk), .CD(n3930), .Q(
        mem_data1[765]) );
  CFD2QXL \mem_data1_reg[766]  ( .D(N10090), .CP(clk), .CD(n3930), .Q(
        mem_data1[766]) );
  CFD2QXL \mem_data1_reg[767]  ( .D(N10091), .CP(clk), .CD(n3930), .Q(
        mem_data1[767]) );
  CFD2QXL \mem_data1_reg[768]  ( .D(N10092), .CP(clk), .CD(n3930), .Q(
        mem_data1[768]) );
  CFD2QXL \mem_data1_reg[769]  ( .D(N10093), .CP(clk), .CD(n3940), .Q(
        mem_data1[769]) );
  CFD2QXL \mem_data1_reg[770]  ( .D(N10094), .CP(clk), .CD(n3930), .Q(
        mem_data1[770]) );
  CFD2QXL \mem_data1_reg[771]  ( .D(N10095), .CP(clk), .CD(n3930), .Q(
        mem_data1[771]) );
  CFD2QXL \mem_data1_reg[772]  ( .D(N10096), .CP(clk), .CD(n3930), .Q(
        mem_data1[772]) );
  CFD2QXL \mem_data1_reg[773]  ( .D(N10097), .CP(clk), .CD(n3930), .Q(
        mem_data1[773]) );
  CFD2QXL \mem_data1_reg[774]  ( .D(N10098), .CP(clk), .CD(n3930), .Q(
        mem_data1[774]) );
  CFD2QXL \mem_data1_reg[775]  ( .D(N10099), .CP(clk), .CD(n3930), .Q(
        mem_data1[775]) );
  CFD2QXL \mem_data1_reg[776]  ( .D(N10100), .CP(clk), .CD(n3930), .Q(
        mem_data1[776]) );
  CFD2QXL \mem_data1_reg[777]  ( .D(N10101), .CP(clk), .CD(n3931), .Q(
        mem_data1[777]) );
  CFD2QXL \mem_data1_reg[778]  ( .D(N10102), .CP(clk), .CD(n3931), .Q(
        mem_data1[778]) );
  CFD2QXL \mem_data1_reg[779]  ( .D(N10103), .CP(clk), .CD(n3931), .Q(
        mem_data1[779]) );
  CFD2QXL \mem_data1_reg[780]  ( .D(N10104), .CP(clk), .CD(n3931), .Q(
        mem_data1[780]) );
  CFD2QXL \mem_data1_reg[781]  ( .D(N10105), .CP(clk), .CD(n3931), .Q(
        mem_data1[781]) );
  CFD2QXL \mem_data1_reg[782]  ( .D(N10106), .CP(clk), .CD(n3931), .Q(
        mem_data1[782]) );
  CFD2QXL \mem_data1_reg[783]  ( .D(N10107), .CP(clk), .CD(n3931), .Q(
        mem_data1[783]) );
  CFD2QXL \mem_data1_reg[784]  ( .D(N10108), .CP(clk), .CD(n3931), .Q(
        mem_data1[784]) );
  CFD2QXL \mem_data1_reg[785]  ( .D(N10109), .CP(clk), .CD(n3931), .Q(
        mem_data1[785]) );
  CFD2QXL \mem_data1_reg[786]  ( .D(N10110), .CP(clk), .CD(n3931), .Q(
        mem_data1[786]) );
  CFD2QXL \mem_data1_reg[787]  ( .D(N10111), .CP(clk), .CD(n3931), .Q(
        mem_data1[787]) );
  CFD2QXL \mem_data1_reg[788]  ( .D(N10112), .CP(clk), .CD(n3931), .Q(
        mem_data1[788]) );
  CFD2QXL \mem_data1_reg[789]  ( .D(N10113), .CP(clk), .CD(n3931), .Q(
        mem_data1[789]) );
  CFD2QXL \mem_data1_reg[790]  ( .D(N10114), .CP(clk), .CD(n3932), .Q(
        mem_data1[790]) );
  CFD2QXL \mem_data1_reg[791]  ( .D(N10115), .CP(clk), .CD(n3932), .Q(
        mem_data1[791]) );
  CFD2QXL \mem_data1_reg[792]  ( .D(N10116), .CP(clk), .CD(n3932), .Q(
        mem_data1[792]) );
  CFD2QXL \mem_data1_reg[793]  ( .D(N10117), .CP(clk), .CD(n3932), .Q(
        mem_data1[793]) );
  CFD2QXL \mem_data1_reg[794]  ( .D(N10118), .CP(clk), .CD(n3932), .Q(
        mem_data1[794]) );
  CFD2QXL \mem_data1_reg[795]  ( .D(N10119), .CP(clk), .CD(n3932), .Q(
        mem_data1[795]) );
  CFD2QXL \mem_data1_reg[796]  ( .D(N10120), .CP(clk), .CD(n3932), .Q(
        mem_data1[796]) );
  CFD2QXL \mem_data1_reg[797]  ( .D(N10121), .CP(clk), .CD(n3932), .Q(
        mem_data1[797]) );
  CFD2QXL \mem_data1_reg[798]  ( .D(N10122), .CP(clk), .CD(n3932), .Q(
        mem_data1[798]) );
  CFD2QXL \mem_data1_reg[799]  ( .D(N10123), .CP(clk), .CD(n3932), .Q(
        mem_data1[799]) );
  CFD2QXL \mem_data1_reg[800]  ( .D(N10124), .CP(clk), .CD(n3932), .Q(
        mem_data1[800]) );
  CFD2QXL \mem_data1_reg[801]  ( .D(N10125), .CP(clk), .CD(n3932), .Q(
        mem_data1[801]) );
  CFD2QXL \mem_data1_reg[802]  ( .D(N10126), .CP(clk), .CD(n3932), .Q(
        mem_data1[802]) );
  CFD2QXL \mem_data1_reg[803]  ( .D(N10127), .CP(clk), .CD(n3933), .Q(
        mem_data1[803]) );
  CFD2QXL \mem_data1_reg[804]  ( .D(N10128), .CP(clk), .CD(n3933), .Q(
        mem_data1[804]) );
  CFD2QXL \mem_data1_reg[805]  ( .D(N10129), .CP(clk), .CD(n3933), .Q(
        mem_data1[805]) );
  CFD2QXL \mem_data1_reg[806]  ( .D(N10130), .CP(clk), .CD(n3933), .Q(
        mem_data1[806]) );
  CFD2QXL \mem_data1_reg[807]  ( .D(N10131), .CP(clk), .CD(n3933), .Q(
        mem_data1[807]) );
  CFD2QXL \mem_data1_reg[808]  ( .D(N10132), .CP(clk), .CD(n3933), .Q(
        mem_data1[808]) );
  CFD2QXL \mem_data1_reg[809]  ( .D(N10133), .CP(clk), .CD(n3933), .Q(
        mem_data1[809]) );
  CFD2QXL \mem_data1_reg[810]  ( .D(N10134), .CP(clk), .CD(n3933), .Q(
        mem_data1[810]) );
  CFD2QXL \mem_data1_reg[811]  ( .D(N10135), .CP(clk), .CD(n3933), .Q(
        mem_data1[811]) );
  CFD2QXL \mem_data1_reg[812]  ( .D(N10136), .CP(clk), .CD(n3933), .Q(
        mem_data1[812]) );
  CFD2QXL \mem_data1_reg[813]  ( .D(N10137), .CP(clk), .CD(n3933), .Q(
        mem_data1[813]) );
  CFD2QXL \mem_data1_reg[814]  ( .D(N10138), .CP(clk), .CD(n3933), .Q(
        mem_data1[814]) );
  CFD2QXL \mem_data1_reg[815]  ( .D(N10139), .CP(clk), .CD(n3933), .Q(
        mem_data1[815]) );
  CFD2QXL \mem_data1_reg[816]  ( .D(N10140), .CP(clk), .CD(n3934), .Q(
        mem_data1[816]) );
  CFD2QXL \mem_data1_reg[817]  ( .D(N10141), .CP(clk), .CD(n3934), .Q(
        mem_data1[817]) );
  CFD2QXL \mem_data1_reg[818]  ( .D(N10142), .CP(clk), .CD(n3934), .Q(
        mem_data1[818]) );
  CFD2QXL \mem_data1_reg[819]  ( .D(N10143), .CP(clk), .CD(n3934), .Q(
        mem_data1[819]) );
  CFD2QXL \mem_data1_reg[820]  ( .D(N10144), .CP(clk), .CD(n3934), .Q(
        mem_data1[820]) );
  CFD2QXL \mem_data1_reg[821]  ( .D(N10145), .CP(clk), .CD(n3934), .Q(
        mem_data1[821]) );
  CFD2QXL \mem_data1_reg[822]  ( .D(N10146), .CP(clk), .CD(n3934), .Q(
        mem_data1[822]) );
  CFD2QXL \mem_data1_reg[823]  ( .D(N10147), .CP(clk), .CD(n3934), .Q(
        mem_data1[823]) );
  CFD2QXL \mem_data1_reg[824]  ( .D(N10148), .CP(clk), .CD(n3934), .Q(
        mem_data1[824]) );
  CFD2QXL \mem_data1_reg[825]  ( .D(N10149), .CP(clk), .CD(n3934), .Q(
        mem_data1[825]) );
  CFD2QXL \mem_data1_reg[826]  ( .D(N10150), .CP(clk), .CD(n3934), .Q(
        mem_data1[826]) );
  CFD2QXL \mem_data1_reg[827]  ( .D(N10151), .CP(clk), .CD(n3934), .Q(
        mem_data1[827]) );
  CFD2QXL \mem_data1_reg[828]  ( .D(N10152), .CP(clk), .CD(n3935), .Q(
        mem_data1[828]) );
  CFD2QXL \mem_data1_reg[829]  ( .D(N10153), .CP(clk), .CD(n3935), .Q(
        mem_data1[829]) );
  CFD2QXL \mem_data1_reg[830]  ( .D(N10154), .CP(clk), .CD(n3935), .Q(
        mem_data1[830]) );
  CFD2QXL \mem_data1_reg[831]  ( .D(N10155), .CP(clk), .CD(n3935), .Q(
        mem_data1[831]) );
  CFD2QXL \mem_data1_reg[832]  ( .D(N10156), .CP(clk), .CD(n3935), .Q(
        mem_data1[832]) );
  CFD2QXL \mem_data1_reg[833]  ( .D(N10157), .CP(clk), .CD(n3935), .Q(
        mem_data1[833]) );
  CFD2QXL \mem_data1_reg[834]  ( .D(N10158), .CP(clk), .CD(n3935), .Q(
        mem_data1[834]) );
  CFD2QXL \mem_data1_reg[835]  ( .D(N10159), .CP(clk), .CD(n3935), .Q(
        mem_data1[835]) );
  CFD2QXL \mem_data1_reg[836]  ( .D(N10160), .CP(clk), .CD(n3935), .Q(
        mem_data1[836]) );
  CFD2QXL \mem_data1_reg[837]  ( .D(N10161), .CP(clk), .CD(n3935), .Q(
        mem_data1[837]) );
  CFD2QXL \mem_data1_reg[838]  ( .D(N10162), .CP(clk), .CD(n3935), .Q(
        mem_data1[838]) );
  CFD2QXL \mem_data1_reg[839]  ( .D(N10163), .CP(clk), .CD(n3935), .Q(
        mem_data1[839]) );
  CFD2QXL \mem_data1_reg[840]  ( .D(N10164), .CP(clk), .CD(n3935), .Q(
        mem_data1[840]) );
  CFD2QXL \mem_data1_reg[841]  ( .D(N10165), .CP(clk), .CD(n3936), .Q(
        mem_data1[841]) );
  CFD2QXL \mem_data1_reg[842]  ( .D(N10166), .CP(clk), .CD(n3936), .Q(
        mem_data1[842]) );
  CFD2QXL \mem_data1_reg[843]  ( .D(N10167), .CP(clk), .CD(n3936), .Q(
        mem_data1[843]) );
  CFD2QXL \mem_data1_reg[844]  ( .D(N10168), .CP(clk), .CD(n3936), .Q(
        mem_data1[844]) );
  CFD2QXL \mem_data1_reg[845]  ( .D(N10169), .CP(clk), .CD(n3936), .Q(
        mem_data1[845]) );
  CFD2QXL \mem_data1_reg[846]  ( .D(N10170), .CP(clk), .CD(n3936), .Q(
        mem_data1[846]) );
  CFD2QXL \mem_data1_reg[847]  ( .D(N10171), .CP(clk), .CD(n3936), .Q(
        mem_data1[847]) );
  CFD2QXL \mem_data1_reg[848]  ( .D(N10172), .CP(clk), .CD(n3936), .Q(
        mem_data1[848]) );
  CFD2QXL \mem_data1_reg[849]  ( .D(N10173), .CP(clk), .CD(n3936), .Q(
        mem_data1[849]) );
  CFD2QXL \mem_data1_reg[850]  ( .D(N10174), .CP(clk), .CD(n3936), .Q(
        mem_data1[850]) );
  CFD2QXL \mem_data1_reg[851]  ( .D(N10175), .CP(clk), .CD(n3936), .Q(
        mem_data1[851]) );
  CFD2QXL \mem_data1_reg[852]  ( .D(N10176), .CP(clk), .CD(n3936), .Q(
        mem_data1[852]) );
  CFD2QXL \mem_data1_reg[853]  ( .D(N10177), .CP(clk), .CD(n3936), .Q(
        mem_data1[853]) );
  CFD2QXL \mem_data1_reg[854]  ( .D(N10178), .CP(clk), .CD(n3937), .Q(
        mem_data1[854]) );
  CFD2QXL \mem_data1_reg[855]  ( .D(N10179), .CP(clk), .CD(n3937), .Q(
        mem_data1[855]) );
  CFD2QXL \mem_data1_reg[856]  ( .D(N10180), .CP(clk), .CD(n3937), .Q(
        mem_data1[856]) );
  CFD2QXL \mem_data1_reg[857]  ( .D(N10181), .CP(clk), .CD(n3937), .Q(
        mem_data1[857]) );
  CFD2QXL \mem_data1_reg[858]  ( .D(N10182), .CP(clk), .CD(n3937), .Q(
        mem_data1[858]) );
  CFD2QXL \mem_data1_reg[859]  ( .D(N10183), .CP(clk), .CD(n3937), .Q(
        mem_data1[859]) );
  CFD2QXL \mem_data1_reg[860]  ( .D(N10184), .CP(clk), .CD(n3937), .Q(
        mem_data1[860]) );
  CFD2QXL \mem_data1_reg[861]  ( .D(N10185), .CP(clk), .CD(n3937), .Q(
        mem_data1[861]) );
  CFD2QXL \mem_data1_reg[862]  ( .D(N10186), .CP(clk), .CD(n3937), .Q(
        mem_data1[862]) );
  CFD2QXL \mem_data1_reg[863]  ( .D(N10187), .CP(clk), .CD(n3937), .Q(
        mem_data1[863]) );
  CFD2QXL \mem_data1_reg[864]  ( .D(N10188), .CP(clk), .CD(n3937), .Q(
        mem_data1[864]) );
  CFD2QXL \mem_data1_reg[865]  ( .D(N10189), .CP(clk), .CD(n3937), .Q(
        mem_data1[865]) );
  CFD2QXL \mem_data1_reg[866]  ( .D(N10190), .CP(clk), .CD(n3937), .Q(
        mem_data1[866]) );
  CFD2QXL \mem_data1_reg[867]  ( .D(N10191), .CP(clk), .CD(n3938), .Q(
        mem_data1[867]) );
  CFD2QXL \mem_data1_reg[868]  ( .D(N10192), .CP(clk), .CD(n3938), .Q(
        mem_data1[868]) );
  CFD2QXL \mem_data1_reg[869]  ( .D(N10193), .CP(clk), .CD(n3938), .Q(
        mem_data1[869]) );
  CFD2QXL \mem_data1_reg[870]  ( .D(N10194), .CP(clk), .CD(n3938), .Q(
        mem_data1[870]) );
  CFD2QXL \mem_data1_reg[871]  ( .D(N10195), .CP(clk), .CD(n3938), .Q(
        mem_data1[871]) );
  CFD2QXL \mem_data1_reg[872]  ( .D(N10196), .CP(clk), .CD(n3938), .Q(
        mem_data1[872]) );
  CFD2QXL \mem_data1_reg[873]  ( .D(N10197), .CP(clk), .CD(n3938), .Q(
        mem_data1[873]) );
  CFD2QXL \mem_data1_reg[874]  ( .D(N10198), .CP(clk), .CD(n3938), .Q(
        mem_data1[874]) );
  CFD2QXL \mem_data1_reg[875]  ( .D(N10199), .CP(clk), .CD(n3938), .Q(
        mem_data1[875]) );
  CFD2QXL \mem_data1_reg[876]  ( .D(N10200), .CP(clk), .CD(n3938), .Q(
        mem_data1[876]) );
  CFD2QXL \mem_data1_reg[877]  ( .D(N10201), .CP(clk), .CD(n3938), .Q(
        mem_data1[877]) );
  CFD2QXL \mem_data1_reg[878]  ( .D(N10202), .CP(clk), .CD(n3938), .Q(
        mem_data1[878]) );
  CFD2QXL \mem_data1_reg[879]  ( .D(N10203), .CP(clk), .CD(n3938), .Q(
        mem_data1[879]) );
  CFD2QXL \mem_data1_reg[880]  ( .D(N10204), .CP(clk), .CD(n3939), .Q(
        mem_data1[880]) );
  CFD2QXL \mem_data1_reg[881]  ( .D(N10205), .CP(clk), .CD(n3939), .Q(
        mem_data1[881]) );
  CFD2QXL \mem_data1_reg[882]  ( .D(N10206), .CP(clk), .CD(n3939), .Q(
        mem_data1[882]) );
  CFD2QXL \mem_data1_reg[883]  ( .D(N10207), .CP(clk), .CD(n3939), .Q(
        mem_data1[883]) );
  CFD2QXL \mem_data1_reg[884]  ( .D(N10208), .CP(clk), .CD(n3939), .Q(
        mem_data1[884]) );
  CFD2QXL \mem_data1_reg[885]  ( .D(N10209), .CP(clk), .CD(n3939), .Q(
        mem_data1[885]) );
  CFD2QXL \mem_data1_reg[886]  ( .D(N10210), .CP(clk), .CD(n3939), .Q(
        mem_data1[886]) );
  CFD2QXL \mem_data1_reg[887]  ( .D(N10211), .CP(clk), .CD(n3939), .Q(
        mem_data1[887]) );
  CFD2QXL \mem_data1_reg[888]  ( .D(N10212), .CP(clk), .CD(n3939), .Q(
        mem_data1[888]) );
  CFD2QXL \mem_data1_reg[889]  ( .D(N10213), .CP(clk), .CD(n3939), .Q(
        mem_data1[889]) );
  CFD2QXL \mem_data1_reg[890]  ( .D(N10214), .CP(clk), .CD(n3939), .Q(
        mem_data1[890]) );
  CFD2QXL \mem_data1_reg[891]  ( .D(N10215), .CP(clk), .CD(n3939), .Q(
        mem_data1[891]) );
  CFD2QXL \mem_data1_reg[892]  ( .D(N10216), .CP(clk), .CD(n3939), .Q(
        mem_data1[892]) );
  CFD2QXL \mem_data1_reg[893]  ( .D(N10217), .CP(clk), .CD(n3940), .Q(
        mem_data1[893]) );
  CFD2QXL \mem_data1_reg[894]  ( .D(N10218), .CP(clk), .CD(n3924), .Q(
        mem_data1[894]) );
  CFD2QXL \mem_data1_reg[895]  ( .D(N10219), .CP(clk), .CD(n3919), .Q(
        mem_data1[895]) );
  CFD2QXL \mem_data1_reg[896]  ( .D(N10220), .CP(clk), .CD(n3919), .Q(
        mem_data1[896]) );
  CFD2QXL \mem_data1_reg[897]  ( .D(N10221), .CP(clk), .CD(n3919), .Q(
        mem_data1[897]) );
  CFD2QXL \mem_data1_reg[898]  ( .D(N10222), .CP(clk), .CD(n3920), .Q(
        mem_data1[898]) );
  CFD2QXL \mem_data1_reg[899]  ( .D(N10223), .CP(clk), .CD(n3920), .Q(
        mem_data1[899]) );
  CFD2QXL \mem_data1_reg[900]  ( .D(N10224), .CP(clk), .CD(n3920), .Q(
        mem_data1[900]) );
  CFD2QXL \mem_data1_reg[901]  ( .D(N10225), .CP(clk), .CD(n3920), .Q(
        mem_data1[901]) );
  CFD2QXL \mem_data1_reg[902]  ( .D(N10226), .CP(clk), .CD(n3920), .Q(
        mem_data1[902]) );
  CFD2QXL \mem_data1_reg[903]  ( .D(N10227), .CP(clk), .CD(n3920), .Q(
        mem_data1[903]) );
  CFD2QXL \mem_data1_reg[904]  ( .D(N10228), .CP(clk), .CD(n3920), .Q(
        mem_data1[904]) );
  CFD2QXL \mem_data1_reg[905]  ( .D(N10229), .CP(clk), .CD(n3920), .Q(
        mem_data1[905]) );
  CFD2QXL \mem_data1_reg[906]  ( .D(N10230), .CP(clk), .CD(n3920), .Q(
        mem_data1[906]) );
  CFD2QXL \mem_data1_reg[907]  ( .D(N10231), .CP(clk), .CD(n3920), .Q(
        mem_data1[907]) );
  CFD2QXL \mem_data1_reg[908]  ( .D(N10232), .CP(clk), .CD(n3920), .Q(
        mem_data1[908]) );
  CFD2QXL \mem_data1_reg[909]  ( .D(N10233), .CP(clk), .CD(n3920), .Q(
        mem_data1[909]) );
  CFD2QXL \mem_data1_reg[910]  ( .D(N10234), .CP(clk), .CD(n3920), .Q(
        mem_data1[910]) );
  CFD2QXL \mem_data1_reg[911]  ( .D(N10235), .CP(clk), .CD(n3921), .Q(
        mem_data1[911]) );
  CFD2QXL \mem_data1_reg[912]  ( .D(N10236), .CP(clk), .CD(n3921), .Q(
        mem_data1[912]) );
  CFD2QXL \mem_data1_reg[913]  ( .D(N10237), .CP(clk), .CD(n3921), .Q(
        mem_data1[913]) );
  CFD2QXL \mem_data1_reg[914]  ( .D(N10238), .CP(clk), .CD(n3921), .Q(
        mem_data1[914]) );
  CFD2QXL \mem_data1_reg[915]  ( .D(N10239), .CP(clk), .CD(n3921), .Q(
        mem_data1[915]) );
  CFD2QXL \mem_data1_reg[916]  ( .D(N10240), .CP(clk), .CD(n3921), .Q(
        mem_data1[916]) );
  CFD2QXL \mem_data1_reg[917]  ( .D(N10241), .CP(clk), .CD(n3921), .Q(
        mem_data1[917]) );
  CFD2QXL \mem_data1_reg[918]  ( .D(N10242), .CP(clk), .CD(n3921), .Q(
        mem_data1[918]) );
  CFD2QXL \mem_data1_reg[919]  ( .D(N10243), .CP(clk), .CD(n3921), .Q(
        mem_data1[919]) );
  CFD2QXL \mem_data1_reg[920]  ( .D(N10244), .CP(clk), .CD(n3921), .Q(
        mem_data1[920]) );
  CFD2QXL \mem_data1_reg[921]  ( .D(N10245), .CP(clk), .CD(n3921), .Q(
        mem_data1[921]) );
  CFD2QXL \mem_data1_reg[922]  ( .D(N10246), .CP(clk), .CD(n3921), .Q(
        mem_data1[922]) );
  CFD2QXL \mem_data1_reg[923]  ( .D(N10247), .CP(clk), .CD(n3921), .Q(
        mem_data1[923]) );
  CFD2QXL \mem_data1_reg[924]  ( .D(N10248), .CP(clk), .CD(n3922), .Q(
        mem_data1[924]) );
  CFD2QXL \mem_data1_reg[925]  ( .D(N10249), .CP(clk), .CD(n3922), .Q(
        mem_data1[925]) );
  CFD2QXL \mem_data1_reg[926]  ( .D(N10250), .CP(clk), .CD(n3922), .Q(
        mem_data1[926]) );
  CFD2QXL \mem_data1_reg[927]  ( .D(N10251), .CP(clk), .CD(n3922), .Q(
        mem_data1[927]) );
  CFD2QXL \mem_data1_reg[928]  ( .D(N10252), .CP(clk), .CD(n3922), .Q(
        mem_data1[928]) );
  CFD2QXL \mem_data1_reg[929]  ( .D(N10253), .CP(clk), .CD(n3922), .Q(
        mem_data1[929]) );
  CFD2QXL \mem_data1_reg[930]  ( .D(N10254), .CP(clk), .CD(n3922), .Q(
        mem_data1[930]) );
  CFD2QXL \mem_data1_reg[931]  ( .D(N10255), .CP(clk), .CD(n3922), .Q(
        mem_data1[931]) );
  CFD2QXL \mem_data1_reg[932]  ( .D(N10256), .CP(clk), .CD(n3922), .Q(
        mem_data1[932]) );
  CFD2QXL \mem_data1_reg[933]  ( .D(N10257), .CP(clk), .CD(n3922), .Q(
        mem_data1[933]) );
  CFD2QXL \mem_data1_reg[934]  ( .D(N10258), .CP(clk), .CD(n3922), .Q(
        mem_data1[934]) );
  CFD2QXL \mem_data1_reg[935]  ( .D(N10259), .CP(clk), .CD(n3922), .Q(
        mem_data1[935]) );
  CFD2QXL \mem_data1_reg[936]  ( .D(N10260), .CP(clk), .CD(n3922), .Q(
        mem_data1[936]) );
  CFD2QXL \mem_data1_reg[937]  ( .D(N10261), .CP(clk), .CD(n3923), .Q(
        mem_data1[937]) );
  CFD2QXL \mem_data1_reg[938]  ( .D(N10262), .CP(clk), .CD(n3923), .Q(
        mem_data1[938]) );
  CFD2QXL \mem_data1_reg[939]  ( .D(N10263), .CP(clk), .CD(n3923), .Q(
        mem_data1[939]) );
  CFD2QXL \mem_data1_reg[940]  ( .D(N10264), .CP(clk), .CD(n3923), .Q(
        mem_data1[940]) );
  CFD2QXL \mem_data1_reg[941]  ( .D(N10265), .CP(clk), .CD(n3923), .Q(
        mem_data1[941]) );
  CFD2QXL \mem_data1_reg[942]  ( .D(N10266), .CP(clk), .CD(n3923), .Q(
        mem_data1[942]) );
  CFD2QXL \mem_data1_reg[943]  ( .D(N10267), .CP(clk), .CD(n3923), .Q(
        mem_data1[943]) );
  CFD2QXL \mem_data1_reg[944]  ( .D(N10268), .CP(clk), .CD(n3923), .Q(
        mem_data1[944]) );
  CFD2QXL \mem_data1_reg[945]  ( .D(N10269), .CP(clk), .CD(n3923), .Q(
        mem_data1[945]) );
  CFD2QXL \mem_data1_reg[946]  ( .D(N10270), .CP(clk), .CD(n3923), .Q(
        mem_data1[946]) );
  CFD2QXL \mem_data1_reg[947]  ( .D(N10271), .CP(clk), .CD(n3923), .Q(
        mem_data1[947]) );
  CFD2QXL \mem_data1_reg[948]  ( .D(N10272), .CP(clk), .CD(n3923), .Q(
        mem_data1[948]) );
  CFD2QXL \mem_data1_reg[949]  ( .D(N10273), .CP(clk), .CD(n3923), .Q(
        mem_data1[949]) );
  CFD2QXL \mem_data1_reg[950]  ( .D(N10274), .CP(clk), .CD(n3924), .Q(
        mem_data1[950]) );
  CFD2QXL \mem_data1_reg[951]  ( .D(N10275), .CP(clk), .CD(n3924), .Q(
        mem_data1[951]) );
  CFD2QXL \mem_data1_reg[952]  ( .D(N10276), .CP(clk), .CD(n3924), .Q(
        mem_data1[952]) );
  CFD2QXL \mem_data1_reg[953]  ( .D(N10277), .CP(clk), .CD(n3924), .Q(
        mem_data1[953]) );
  CFD2QXL \mem_data1_reg[954]  ( .D(N10278), .CP(clk), .CD(n3924), .Q(
        mem_data1[954]) );
  CFD2QXL \mem_data1_reg[955]  ( .D(N10279), .CP(clk), .CD(n3924), .Q(
        mem_data1[955]) );
  CFD2QXL \mem_data1_reg[956]  ( .D(N10280), .CP(clk), .CD(n3924), .Q(
        mem_data1[956]) );
  CFD2QXL \mem_data1_reg[958]  ( .D(N10282), .CP(clk), .CD(n3924), .Q(
        mem_data1[958]) );
  CFD2QXL \mem_data1_reg[959]  ( .D(N10283), .CP(clk), .CD(n3924), .Q(
        mem_data1[959]) );
  CFD2QXL \mem_data1_reg[960]  ( .D(N10284), .CP(clk), .CD(n3924), .Q(
        mem_data1[960]) );
  CFD2QXL \mem_data1_reg[961]  ( .D(N10285), .CP(clk), .CD(n3924), .Q(
        mem_data1[961]) );
  CFD2QXL \mem_data1_reg[962]  ( .D(N10286), .CP(clk), .CD(n3925), .Q(
        mem_data1[962]) );
  CFD2QXL \mem_data1_reg[963]  ( .D(N10287), .CP(clk), .CD(n3925), .Q(
        mem_data1[963]) );
  CFD2QXL \mem_data1_reg[964]  ( .D(N10288), .CP(clk), .CD(n3925), .Q(
        mem_data1[964]) );
  CFD2QXL \mem_data1_reg[965]  ( .D(N10289), .CP(clk), .CD(n3925), .Q(
        mem_data1[965]) );
  CFD2QXL \mem_data1_reg[966]  ( .D(N10290), .CP(clk), .CD(n3925), .Q(
        mem_data1[966]) );
  CFD2QXL \mem_data1_reg[967]  ( .D(N10291), .CP(clk), .CD(n3925), .Q(
        mem_data1[967]) );
  CFD2QXL \mem_data1_reg[968]  ( .D(N10292), .CP(clk), .CD(n3925), .Q(
        mem_data1[968]) );
  CFD2QXL \mem_data1_reg[969]  ( .D(N10293), .CP(clk), .CD(n3925), .Q(
        mem_data1[969]) );
  CFD2QXL \mem_data1_reg[970]  ( .D(N10294), .CP(clk), .CD(n3925), .Q(
        mem_data1[970]) );
  CFD2QXL \mem_data1_reg[971]  ( .D(N10295), .CP(clk), .CD(n3925), .Q(
        mem_data1[971]) );
  CFD2QXL \mem_data1_reg[972]  ( .D(N10296), .CP(clk), .CD(n3925), .Q(
        mem_data1[972]) );
  CFD2QXL \mem_data1_reg[973]  ( .D(N10297), .CP(clk), .CD(n3925), .Q(
        mem_data1[973]) );
  CFD2QXL \mem_data1_reg[974]  ( .D(N10298), .CP(clk), .CD(n3925), .Q(
        mem_data1[974]) );
  CFD2QXL \mem_data1_reg[975]  ( .D(N10299), .CP(clk), .CD(n3926), .Q(
        mem_data1[975]) );
  CFD2QXL \mem_data1_reg[976]  ( .D(N10300), .CP(clk), .CD(n3926), .Q(
        mem_data1[976]) );
  CFD2QXL \mem_data1_reg[977]  ( .D(N10301), .CP(clk), .CD(n3926), .Q(
        mem_data1[977]) );
  CFD2QXL \mem_data1_reg[978]  ( .D(N10302), .CP(clk), .CD(n3926), .Q(
        mem_data1[978]) );
  CFD2QXL \mem_data1_reg[979]  ( .D(N10303), .CP(clk), .CD(n3926), .Q(
        mem_data1[979]) );
  CFD2QXL \mem_data1_reg[980]  ( .D(N10304), .CP(clk), .CD(n3926), .Q(
        mem_data1[980]) );
  CFD2QXL \mem_data1_reg[981]  ( .D(N10305), .CP(clk), .CD(n3926), .Q(
        mem_data1[981]) );
  CFD2QXL \mem_data1_reg[982]  ( .D(N10306), .CP(clk), .CD(n3926), .Q(
        mem_data1[982]) );
  CFD2QXL \mem_data1_reg[983]  ( .D(N10307), .CP(clk), .CD(n3926), .Q(
        mem_data1[983]) );
  CFD2QXL \mem_data1_reg[984]  ( .D(N10308), .CP(clk), .CD(n3926), .Q(
        mem_data1[984]) );
  CFD2QXL \mem_data1_reg[985]  ( .D(N10309), .CP(clk), .CD(n3926), .Q(
        mem_data1[985]) );
  CFD2QXL \mem_data1_reg[986]  ( .D(N10310), .CP(clk), .CD(n3926), .Q(
        mem_data1[986]) );
  CFD2QXL \mem_data1_reg[987]  ( .D(N10311), .CP(clk), .CD(n3926), .Q(
        mem_data1[987]) );
  CFD2QXL \mem_data1_reg[988]  ( .D(N10312), .CP(clk), .CD(n3927), .Q(
        mem_data1[988]) );
  CFD2QXL \mem_data1_reg[989]  ( .D(N10313), .CP(clk), .CD(n3927), .Q(
        mem_data1[989]) );
  CFD2QXL \mem_data1_reg[990]  ( .D(N10314), .CP(clk), .CD(n3927), .Q(
        mem_data1[990]) );
  CFD2QXL \mem_data1_reg[991]  ( .D(N10315), .CP(clk), .CD(n3927), .Q(
        mem_data1[991]) );
  CFD2QXL \mem_data1_reg[992]  ( .D(N10316), .CP(clk), .CD(n3927), .Q(
        mem_data1[992]) );
  CFD2QXL \mem_data1_reg[993]  ( .D(N10317), .CP(clk), .CD(n3927), .Q(
        mem_data1[993]) );
  CFD2QXL \mem_data1_reg[994]  ( .D(N10318), .CP(clk), .CD(n3927), .Q(
        mem_data1[994]) );
  CFD2QXL \mem_data1_reg[995]  ( .D(N10319), .CP(clk), .CD(n3927), .Q(
        mem_data1[995]) );
  CFD2QXL \mem_data1_reg[996]  ( .D(N10320), .CP(clk), .CD(n3927), .Q(
        mem_data1[996]) );
  CFD2QXL \mem_data1_reg[997]  ( .D(N10321), .CP(clk), .CD(n3927), .Q(
        mem_data1[997]) );
  CFD2QXL \mem_data1_reg[998]  ( .D(N10322), .CP(clk), .CD(n3927), .Q(
        mem_data1[998]) );
  CFD2QXL \mem_data1_reg[999]  ( .D(N10323), .CP(clk), .CD(n3927), .Q(
        mem_data1[999]) );
  CFD2QXL \mem_data1_reg[1000]  ( .D(N10324), .CP(clk), .CD(n3927), .Q(
        mem_data1[1000]) );
  CFD2QXL \mem_data1_reg[1001]  ( .D(N10325), .CP(clk), .CD(n3928), .Q(
        mem_data1[1001]) );
  CFD2QXL \mem_data1_reg[1002]  ( .D(N10326), .CP(clk), .CD(n3928), .Q(
        mem_data1[1002]) );
  CFD2QXL \mem_data1_reg[1003]  ( .D(N10327), .CP(clk), .CD(n3928), .Q(
        mem_data1[1003]) );
  CFD2QXL \mem_data1_reg[1004]  ( .D(N10328), .CP(clk), .CD(n3928), .Q(
        mem_data1[1004]) );
  CFD2QXL \mem_data1_reg[1005]  ( .D(N10329), .CP(clk), .CD(n3928), .Q(
        mem_data1[1005]) );
  CFD2QXL \mem_data1_reg[1006]  ( .D(N10330), .CP(clk), .CD(n3928), .Q(
        mem_data1[1006]) );
  CFD2QXL \mem_data1_reg[1007]  ( .D(N10331), .CP(clk), .CD(n3928), .Q(
        mem_data1[1007]) );
  CFD2QXL \mem_data1_reg[1008]  ( .D(N10332), .CP(clk), .CD(n3928), .Q(
        mem_data1[1008]) );
  CFD2QXL \mem_data1_reg[1009]  ( .D(N10333), .CP(clk), .CD(n3928), .Q(
        mem_data1[1009]) );
  CFD2QXL \mem_data1_reg[1010]  ( .D(N10334), .CP(clk), .CD(n3928), .Q(
        mem_data1[1010]) );
  CFD2QXL \mem_data1_reg[1011]  ( .D(N10335), .CP(clk), .CD(n3928), .Q(
        mem_data1[1011]) );
  CFD2QXL \mem_data1_reg[1012]  ( .D(N10336), .CP(clk), .CD(n3928), .Q(
        mem_data1[1012]) );
  CFD2QXL \mem_data1_reg[1013]  ( .D(N10337), .CP(clk), .CD(n3928), .Q(
        mem_data1[1013]) );
  CFD2QXL \mem_data1_reg[1014]  ( .D(N10338), .CP(clk), .CD(n3929), .Q(
        mem_data1[1014]) );
  CFD2QXL \mem_data1_reg[1015]  ( .D(N10339), .CP(clk), .CD(n3929), .Q(
        mem_data1[1015]) );
  CFD2QXL \mem_data1_reg[1016]  ( .D(N10340), .CP(clk), .CD(n3929), .Q(
        mem_data1[1016]) );
  CFD2QXL \mem_data1_reg[1017]  ( .D(N10341), .CP(clk), .CD(n3929), .Q(
        mem_data1[1017]) );
  CFD2QXL \mem_data1_reg[1018]  ( .D(N10342), .CP(clk), .CD(n3929), .Q(
        mem_data1[1018]) );
  CFD2QXL \mem_data1_reg[1019]  ( .D(N10343), .CP(clk), .CD(n3929), .Q(
        mem_data1[1019]) );
  CFD2QXL \mem_data1_reg[1020]  ( .D(N10344), .CP(clk), .CD(n3929), .Q(
        mem_data1[1020]) );
  CFD2QXL \mem_data1_reg[1021]  ( .D(N10345), .CP(clk), .CD(n3929), .Q(
        mem_data1[1021]) );
  CFD2QXL \mem_data1_reg[319]  ( .D(N9643), .CP(clk), .CD(n3978), .Q(
        mem_data1[319]) );
  CFD2QXL \mem_data1_reg[418]  ( .D(N9742), .CP(clk), .CD(n3965), .Q(
        mem_data1[418]) );
  CFD2QXL \mem_data1_reg[422]  ( .D(N9746), .CP(clk), .CD(n3965), .Q(
        mem_data1[422]) );
  CFD2QXL \mem_data1_reg[447]  ( .D(N9771), .CP(clk), .CD(n3967), .Q(
        mem_data1[447]) );
  CFD2QXL \mem_data1_reg[14]  ( .D(N9338), .CP(clk), .CD(n3954), .Q(
        mem_data1[14]) );
  CFD2QXL \mem_data1_reg[4]  ( .D(N9328), .CP(clk), .CD(n3954), .Q(
        mem_data1[4]) );
  CFD2QXL \mem_data1_reg[11]  ( .D(N9335), .CP(clk), .CD(n3954), .Q(
        mem_data1[11]) );
  CFD2QXL \mem_data1_reg[12]  ( .D(N9336), .CP(clk), .CD(n3954), .Q(
        mem_data1[12]) );
  CFD2QXL \mem_data1_reg[13]  ( .D(N9337), .CP(clk), .CD(n3954), .Q(
        mem_data1[13]) );
  CFD2QXL \mem_data1_reg[10]  ( .D(N9334), .CP(clk), .CD(n3954), .Q(
        mem_data1[10]) );
  CFD2QXL \mem_data1_reg[1]  ( .D(N9325), .CP(clk), .CD(n3953), .Q(
        mem_data1[1]) );
  CFD2QXL \mem_data1_reg[3]  ( .D(N9327), .CP(clk), .CD(n3954), .Q(
        mem_data1[3]) );
  CFD2QXL \mem_data1_reg[5]  ( .D(N9329), .CP(clk), .CD(n3954), .Q(
        mem_data1[5]) );
  CFD2QXL \mem_data1_reg[6]  ( .D(N9330), .CP(clk), .CD(n3954), .Q(
        mem_data1[6]) );
  CFD2QXL \mem_data1_reg[7]  ( .D(N9331), .CP(clk), .CD(n3954), .Q(
        mem_data1[7]) );
  CFD2QXL \mem_data1_reg[8]  ( .D(N9332), .CP(clk), .CD(n3954), .Q(
        mem_data1[8]) );
  CFD2QXL \mem_data1_reg[9]  ( .D(N9333), .CP(clk), .CD(n3954), .Q(
        mem_data1[9]) );
  CFD2QXL \mem_data1_reg[2]  ( .D(N9326), .CP(clk), .CD(n3954), .Q(
        mem_data1[2]) );
  CFD2QXL \mem_data1_reg[253]  ( .D(N9577), .CP(clk), .CD(n3973), .Q(
        mem_data1[253]) );
  CFD2QXL \mem_data1_reg[291]  ( .D(N9615), .CP(clk), .CD(n3976), .Q(
        mem_data1[291]) );
  CFD2QXL \mem_data1_reg[297]  ( .D(N9621), .CP(clk), .CD(n3976), .Q(
        mem_data1[297]) );
  CFD2QXL \mem_data1_reg[298]  ( .D(N9622), .CP(clk), .CD(n3976), .Q(
        mem_data1[298]) );
  CFD2QXL \mem_data1_reg[300]  ( .D(N9624), .CP(clk), .CD(n3977), .Q(
        mem_data1[300]) );
  CFD2QXL \mem_data1_reg[417]  ( .D(N9741), .CP(clk), .CD(n3965), .Q(
        mem_data1[417]) );
  CFD2QXL \mem_data1_reg[419]  ( .D(N9743), .CP(clk), .CD(n3965), .Q(
        mem_data1[419]) );
  CFD2QXL \mem_data1_reg[436]  ( .D(N9760), .CP(clk), .CD(n3966), .Q(
        mem_data1[436]) );
  CFD2QXL \mem_data1_reg[437]  ( .D(N9761), .CP(clk), .CD(n3966), .Q(
        mem_data1[437]) );
  CFD2QXL \mem_data1_reg[441]  ( .D(N9765), .CP(clk), .CD(n3967), .Q(
        mem_data1[441]) );
  CFD2QXL \mem_data1_reg[442]  ( .D(N9766), .CP(clk), .CD(n3967), .Q(
        mem_data1[442]) );
  CFD2QXL \mem_data1_reg[443]  ( .D(N9767), .CP(clk), .CD(n3967), .Q(
        mem_data1[443]) );
  CFD2QXL \mem_data1_reg[444]  ( .D(N9768), .CP(clk), .CD(n3967), .Q(
        mem_data1[444]) );
  CFD2QXL \mem_data1_reg[446]  ( .D(N9770), .CP(clk), .CD(n3967), .Q(
        mem_data1[446]) );
  CFD2QXL \mem_data1_reg[485]  ( .D(N9809), .CP(clk), .CD(n3970), .Q(
        mem_data1[485]) );
  CFD2QXL \mem_data1_reg[255]  ( .D(N9579), .CP(clk), .CD(n3973), .Q(
        mem_data1[255]) );
  CFD2QXL \mem_data1_reg[383]  ( .D(N9707), .CP(clk), .CD(n3962), .Q(
        mem_data1[383]) );
  CFD2QXL \mem_data1_reg[487]  ( .D(N9811), .CP(clk), .CD(n3970), .Q(
        mem_data1[487]) );
  CFD2QXL \datain0_reg[31]  ( .D(datain[31]), .CP(clk), .CD(n3950), .Q(
        datain0[31]) );
  CFD2QXL \datain0_reg[30]  ( .D(datain[30]), .CP(clk), .CD(n3950), .Q(
        datain0[30]) );
  CFD2QXL \datain0_reg[29]  ( .D(datain[29]), .CP(clk), .CD(n3950), .Q(
        datain0[29]) );
  CFD2QXL \datain0_reg[28]  ( .D(datain[28]), .CP(clk), .CD(n3950), .Q(
        datain0[28]) );
  CFD2QXL \datain0_reg[27]  ( .D(datain[27]), .CP(clk), .CD(n3950), .Q(
        datain0[27]) );
  CFD2QXL \datain0_reg[26]  ( .D(datain[26]), .CP(clk), .CD(n3951), .Q(
        datain0[26]) );
  CFD2QXL \datain0_reg[25]  ( .D(datain[25]), .CP(clk), .CD(n3951), .Q(
        datain0[25]) );
  CFD2QXL \datain0_reg[8]  ( .D(datain[8]), .CP(clk), .CD(n3952), .Q(
        datain0[8]) );
  CFD2QXL \datain0_reg[6]  ( .D(datain[6]), .CP(clk), .CD(n3952), .Q(
        datain0[6]) );
  CFD2QXL \datain0_reg[5]  ( .D(datain[5]), .CP(clk), .CD(n3952), .Q(
        datain0[5]) );
  CFD2QXL \datain0_reg[4]  ( .D(datain[4]), .CP(clk), .CD(n3952), .Q(
        datain0[4]) );
  CFD2QXL \datain0_reg[3]  ( .D(datain[3]), .CP(clk), .CD(n3952), .Q(
        datain0[3]) );
  CFD2QXL \datain0_reg[2]  ( .D(datain[2]), .CP(clk), .CD(n3952), .Q(
        datain0[2]) );
  CFD2QXL \datain0_reg[1]  ( .D(datain[1]), .CP(clk), .CD(n3952), .Q(
        datain0[1]) );
  CFD2QXL \datain0_reg[0]  ( .D(datain[0]), .CP(clk), .CD(n3953), .Q(
        datain0[0]) );
  CFD2QXL \wr_ptr_reg[2]  ( .D(N10350), .CP(clk), .CD(n3953), .Q(N2068) );
  CFD2QXL \datain0_reg[24]  ( .D(datain[24]), .CP(clk), .CD(n3951), .Q(
        datain0[24]) );
  CFD2QXL \datain0_reg[23]  ( .D(datain[23]), .CP(clk), .CD(n3951), .Q(
        datain0[23]) );
  CFD2QXL \datain0_reg[22]  ( .D(datain[22]), .CP(clk), .CD(n3951), .Q(
        datain0[22]) );
  CFD2QXL \datain0_reg[21]  ( .D(datain[21]), .CP(clk), .CD(n3951), .Q(
        datain0[21]) );
  CFD2QXL \datain0_reg[20]  ( .D(datain[20]), .CP(clk), .CD(n3951), .Q(
        datain0[20]) );
  CFD2QXL \datain0_reg[19]  ( .D(datain[19]), .CP(clk), .CD(n3951), .Q(
        datain0[19]) );
  CFD2QXL \datain0_reg[18]  ( .D(datain[18]), .CP(clk), .CD(n3951), .Q(
        datain0[18]) );
  CFD2QXL \datain0_reg[17]  ( .D(datain[17]), .CP(clk), .CD(n3951), .Q(
        datain0[17]) );
  CFD2QXL \datain0_reg[16]  ( .D(datain[16]), .CP(clk), .CD(n3951), .Q(
        datain0[16]) );
  CFD2QXL \datain0_reg[15]  ( .D(datain[15]), .CP(clk), .CD(n3951), .Q(
        datain0[15]) );
  CFD2QXL \datain0_reg[14]  ( .D(datain[14]), .CP(clk), .CD(n3951), .Q(
        datain0[14]) );
  CFD2QXL \datain0_reg[13]  ( .D(datain[13]), .CP(clk), .CD(n3952), .Q(
        datain0[13]) );
  CFD2QXL \datain0_reg[12]  ( .D(datain[12]), .CP(clk), .CD(n3952), .Q(
        datain0[12]) );
  CFD2QXL \datain0_reg[11]  ( .D(datain[11]), .CP(clk), .CD(n3952), .Q(
        datain0[11]) );
  CFD2QXL \datain0_reg[10]  ( .D(datain[10]), .CP(clk), .CD(n3952), .Q(
        datain0[10]) );
  CFD2QXL \datain0_reg[9]  ( .D(datain[9]), .CP(clk), .CD(n3952), .Q(
        datain0[9]) );
  CFD2QXL \datain0_reg[7]  ( .D(datain[7]), .CP(clk), .CD(n3952), .Q(
        datain0[7]) );
  CFD2QXL \lenin01_reg[3]  ( .D(n3533), .CP(clk), .CD(n3929), .Q(lenout[3]) );
  CFD2XL pushout_reg_reg ( .D(N10358), .CP(clk), .CD(n3899), .Q(pushout), .QN(
        n52) );
  CFD2QX1 \lenin0_reg[0]  ( .D(reqlen[0]), .CP(clk), .CD(n3950), .Q(lenin0[0])
         );
  CFD2QX1 \wr_ptr_reg[1]  ( .D(N10349), .CP(clk), .CD(n3953), .Q(N2067) );
  CFD4QXL \wr_ptr_reg[8]  ( .D(N10356), .CP(clk), .SD(n3981), .Q(wr_ptr[8]) );
  CFD2XL \dataout_reg1_reg[14]  ( .D(n3173), .CP(clk), .CD(n4415), .QN(n37) );
  CFD2XL \dataout_reg1_reg[13]  ( .D(n3174), .CP(clk), .CD(n4415), .QN(n38) );
  CFD2XL \dataout_reg1_reg[12]  ( .D(n3175), .CP(clk), .CD(n4415), .QN(n39) );
  CFD2XL \dataout_reg1_reg[11]  ( .D(n3176), .CP(clk), .CD(n4415), .QN(n40) );
  CFD2XL \dataout_reg1_reg[10]  ( .D(n3177), .CP(clk), .CD(n4415), .QN(n41) );
  CFD2XL \dataout_reg1_reg[9]  ( .D(n3178), .CP(clk), .CD(n4415), .QN(n42) );
  CFD2XL \dataout_reg1_reg[8]  ( .D(n3179), .CP(clk), .CD(n4415), .QN(n43) );
  CFD2XL \dataout_reg1_reg[7]  ( .D(n3180), .CP(clk), .CD(n4415), .QN(n44) );
  CFD2XL \dataout_reg1_reg[6]  ( .D(n3181), .CP(clk), .CD(n4415), .QN(n45) );
  CFD2XL \dataout_reg1_reg[5]  ( .D(n3182), .CP(clk), .CD(n4415), .QN(n46) );
  CFD2XL \dataout_reg1_reg[4]  ( .D(n3183), .CP(clk), .CD(n4415), .QN(n47) );
  CFD2XL \dataout_reg1_reg[3]  ( .D(n3184), .CP(clk), .CD(n4415), .QN(n48) );
  CFD2XL \dataout_reg1_reg[2]  ( .D(n3185), .CP(clk), .CD(n4415), .QN(n49) );
  CFD2XL \dataout_reg1_reg[1]  ( .D(n3186), .CP(clk), .CD(n4415), .QN(n50) );
  CFD2XL \dataout_reg1_reg[0]  ( .D(n3187), .CP(clk), .CD(n4415), .QN(n51) );
  CFD4QXL \wr_ptr_reg[6]  ( .D(N10354), .CP(clk), .SD(n4415), .Q(wr_ptr[6]) );
  CFD2XL \lenin01_reg[1]  ( .D(n3223), .CP(clk), .CD(n4415), .Q(lenout[1]), 
        .QN(n4440) );
  CFD2QXL \lenin0_reg[1]  ( .D(reqlen[1]), .CP(clk), .CD(n3955), .Q(lenin0[1])
         );
  CFD4QX2 \wr_ptr_reg[9]  ( .D(N10357), .CP(clk), .SD(n3981), .Q(wr_ptr[9]) );
  CFD2QX1 \wr_ptr_reg[0]  ( .D(N10348), .CP(clk), .CD(n3953), .Q(N2066) );
  CFD4QXL \wr_ptr_reg[5]  ( .D(N10353), .CP(clk), .SD(n3981), .Q(wr_ptr[5]) );
  CFD2QXL pushin0_reg ( .D(pushin), .CP(clk), .CD(n3953), .Q(pushin0) );
  CFD2QXL reqin0_reg ( .D(reqin), .CP(clk), .CD(n3953), .Q(reqin0) );
  CFD2QXL \lenin0_reg[3]  ( .D(reqlen[3]), .CP(clk), .CD(n3899), .Q(lenin0[3])
         );
  CFD4QXL \wr_ptr_reg[7]  ( .D(N10355), .CP(clk), .SD(n3981), .Q(wr_ptr[7]) );
  CIVDX2 U5222 ( .A(N2067), .Z0(n3188), .Z1(n3189) );
  CIVDX2 U5223 ( .A(N2067), .Z0(n3190), .Z1(n3191) );
  CIVDX2 U5224 ( .A(N2067), .Z0(n3192), .Z1(n3193) );
  CIVDX2 U5225 ( .A(N2067), .Z0(n3194), .Z1(n3195) );
  CIVX2 U5226 ( .A(wr_ptr[5]), .Z(n3196) );
  CIVX1 U5227 ( .A(wr_ptr[5]), .Z(n3197) );
  CIVXL U5228 ( .A(wr_ptr[5]), .Z(n3198) );
  CIVDX4 U5229 ( .A(n3196), .Z0(n3199), .Z1(n3200) );
  CIVDX1 U5230 ( .A(n3196), .Z0(n3201), .Z1(n3202) );
  CIVDX1 U5231 ( .A(n3196), .Z0(n3203), .Z1(n3204) );
  CIVDX1 U5232 ( .A(n3197), .Z0(n3205), .Z1(n3206) );
  CIVDX1 U5233 ( .A(n3197), .Z0(n3207), .Z1(n3208) );
  CIVDX1 U5234 ( .A(n3197), .Z0(n3209), .Z1(n3210) );
  CIVDX1 U5235 ( .A(n3198), .Z0(n3211), .Z1(n3212) );
  CIVDX1 U5236 ( .A(n3198), .Z0(n3213), .Z1(n3214) );
  CIVDX1 U5237 ( .A(n3198), .Z0(n3215), .Z1(n3216) );
  CIVX2 U5238 ( .A(N2066), .Z(n4436) );
  COR4X1 U5239 ( .A(lenin0[1]), .B(n4294), .C(n3533), .D(lenin0[2]), .Z(n3171)
         );
  CNIVX1 U5240 ( .A(n4302), .Z(n4299) );
  CNIVX1 U5241 ( .A(n4304), .Z(n4295) );
  CNIVX1 U5242 ( .A(n4378), .Z(n4384) );
  CNIVX1 U5243 ( .A(n4378), .Z(n4380) );
  CNIVX1 U5244 ( .A(n4378), .Z(n4382) );
  CNIVX1 U5245 ( .A(n4377), .Z(n4379) );
  CNIVX1 U5246 ( .A(n74), .Z(n3640) );
  CIVX2 U5247 ( .A(mem_data1[434]), .Z(n3241) );
  CNR4X1 U5248 ( .A(n3640), .B(n3217), .C(n3570), .D(n3606), .Z(n75) );
  CNIVX1 U5249 ( .A(n3769), .Z(n4383) );
  CNIVX1 U5250 ( .A(n4377), .Z(n4381) );
  CNIVX1 U5251 ( .A(n4302), .Z(n4300) );
  CNIVX1 U5252 ( .A(n4303), .Z(n4296) );
  CNIVX1 U5253 ( .A(n4303), .Z(n4298) );
  CNIVX1 U5254 ( .A(n4303), .Z(n4297) );
  CAN2X1 U5255 ( .A(n3170), .B(n3222), .Z(n3217) );
  CNIVX1 U5256 ( .A(N2069), .Z(n3754) );
  CIVX2 U5257 ( .A(wr_ptr[8]), .Z(n4390) );
  CIVDX1 U5258 ( .A(wr_ptr[6]), .Z0(n3720), .Z1(n3721) );
  CMX2X1 U5259 ( .A0(n4642), .A1(n4644), .S(n4227), .Z(n3219) );
  COR2X1 U5260 ( .A(n4434), .B(n4435), .Z(n3220) );
  COR2X1 U5261 ( .A(n3171), .B(n3220), .Z(n3221) );
  CNIVX1 U5262 ( .A(n3756), .Z(n3757) );
  CAN2X1 U5263 ( .A(reqin0), .B(pushin0), .Z(n3222) );
  CNIVX1 U5264 ( .A(n3750), .Z(n3223) );
  CNIVX1 U5265 ( .A(n51), .Z(n3224) );
  CNIVX1 U5266 ( .A(n50), .Z(n3225) );
  CNIVX1 U5267 ( .A(n49), .Z(n3226) );
  CNIVX1 U5268 ( .A(n48), .Z(n3227) );
  CNIVX1 U5269 ( .A(n47), .Z(n3228) );
  CNIVX1 U5270 ( .A(n46), .Z(n3229) );
  CNIVX1 U5271 ( .A(n45), .Z(n3230) );
  CNIVX1 U5272 ( .A(n44), .Z(n3231) );
  CNIVX1 U5273 ( .A(n43), .Z(n3232) );
  CNIVX1 U5274 ( .A(n42), .Z(n3233) );
  CNIVX1 U5275 ( .A(n41), .Z(n3234) );
  CNIVX1 U5276 ( .A(n40), .Z(n3235) );
  CNIVX1 U5277 ( .A(n39), .Z(n3236) );
  CNIVX1 U5278 ( .A(n38), .Z(n3237) );
  CNIVX1 U5279 ( .A(n37), .Z(n3238) );
  CMXI2XL U5280 ( .A0(n4718), .A1(n4720), .S(n3763), .Z(n4704) );
  CIVXL U5281 ( .A(n4720), .Z(n3701) );
  CENX1 U5282 ( .A(n3239), .B(mem_data1[155]), .Z(N8124) );
  COR2X1 U5283 ( .A(n3829), .B(n5170), .Z(n3239) );
  CNR2X1 U5284 ( .A(n3741), .B(n3757), .Z(n3240) );
  CMXI2XL U5285 ( .A0(n5022), .A1(n4994), .S(n4219), .Z(n5052) );
  CMXI2X1 U5286 ( .A0(n13848), .A1(n13871), .S(n3533), .Z(N8711) );
  CENX1 U5287 ( .A(N452), .B(n3241), .Z(N7845) );
  CANR2XL U5288 ( .A(N2345), .B(n3586), .C(n3621), .D(N8010), .Z(n1297) );
  CMX2XL U5289 ( .A0(N8010), .A1(N8009), .S(n4240), .Z(n10184) );
  CMX2XL U5290 ( .A0(N8011), .A1(N8010), .S(n4242), .Z(n10181) );
  CMXI2X1 U5291 ( .A0(n4938), .A1(n4920), .S(n4217), .Z(n4963) );
  CMXI2XL U5292 ( .A0(n4928), .A1(n4919), .S(n3188), .Z(n4938) );
  CNIVXL U5293 ( .A(n4437), .Z(n3247) );
  CNIVXL U5294 ( .A(n4437), .Z(n3246) );
  CNIVXL U5295 ( .A(n4437), .Z(n4214) );
  CNR2XL U5296 ( .A(n6044), .B(n4215), .Z(n6065) );
  CNR2XL U5297 ( .A(n5480), .B(n4218), .Z(n5501) );
  COR2X1 U5298 ( .A(N3107), .B(\r349/carry [7]), .Z(\r349/carry [8]) );
  CENX1 U5299 ( .A(N3107), .B(\r349/carry [7]), .Z(N6229) );
  CND2X1 U5300 ( .A(n6046), .B(n4406), .Z(n6052) );
  CND2X1 U5301 ( .A(n6051), .B(n4408), .Z(n6057) );
  CIVXL U5302 ( .A(n3219), .Z(n3242) );
  CND2X1 U5303 ( .A(n3830), .B(n3243), .Z(n3244) );
  CND2XL U5304 ( .A(n3851), .B(\r347/carry [7]), .Z(n3245) );
  CND2X1 U5305 ( .A(n3244), .B(n3245), .Z(N3107) );
  CIVXL U5306 ( .A(\r347/carry [7]), .Z(n3243) );
  CAN2XL U5307 ( .A(N2066), .B(n4293), .Z(\r347/carry [1]) );
  CIVX2 U5308 ( .A(n4301), .Z(n4293) );
  CMXI2X1 U5309 ( .A0(n15725), .A1(n12712), .S(n3271), .Z(N9287) );
  CMXI2X1 U5310 ( .A0(n15723), .A1(n12710), .S(n3271), .Z(N9286) );
  CMXI2XL U5311 ( .A0(n12712), .A1(n12720), .S(n3532), .Z(N9295) );
  CMXI2XL U5312 ( .A0(n12710), .A1(n12719), .S(n3394), .Z(N9294) );
  CNR2XL U5313 ( .A(n3508), .B(n9643), .Z(N6176) );
  CNR2XL U5314 ( .A(n3450), .B(n9641), .Z(N6174) );
  CNR2XL U5315 ( .A(n3270), .B(n9642), .Z(N6175) );
  CNR2XL U5316 ( .A(n3270), .B(n9644), .Z(N6177) );
  CNR2X1 U5317 ( .A(n4718), .B(n3759), .Z(n4795) );
  CND2X1 U5318 ( .A(n4886), .B(n3735), .Z(n6155) );
  CND2X1 U5319 ( .A(n4887), .B(n3738), .Z(n6182) );
  CND2X1 U5320 ( .A(n4885), .B(n3733), .Z(n6125) );
  CND2X1 U5321 ( .A(n5255), .B(n3728), .Z(n5356) );
  CND2IX1 U5322 ( .B(n5198), .A(n3723), .Z(n5300) );
  CNR2XL U5323 ( .A(n4749), .B(n3760), .Z(n4778) );
  CNIVX1 U5324 ( .A(n79), .Z(n3606) );
  CNIVX1 U5325 ( .A(n73), .Z(n3570) );
  CMX2X1 U5326 ( .A0(N7279), .A1(N7278), .S(n3880), .Z(n15690) );
  CMX2XL U5327 ( .A0(N7281), .A1(N7280), .S(n3863), .Z(n15689) );
  CIVX4 U5328 ( .A(n3896), .Z(n4437) );
  CNR2XL U5329 ( .A(n4216), .B(n4929), .Z(n4951) );
  CNIVXL U5330 ( .A(n79), .Z(n3636) );
  CNIVXL U5331 ( .A(n79), .Z(n3610) );
  CNIVXL U5332 ( .A(n79), .Z(n3612) );
  CNIVXL U5333 ( .A(n73), .Z(n3576) );
  CNIVXL U5334 ( .A(n73), .Z(n3603) );
  CNIVXL U5335 ( .A(n73), .Z(n3573) );
  CNIVXL U5336 ( .A(n73), .Z(n3584) );
  CNIVXL U5337 ( .A(n79), .Z(n3633) );
  CNIVXL U5338 ( .A(n79), .Z(n3620) );
  CNIVXL U5339 ( .A(n79), .Z(n3618) );
  CNIVXL U5340 ( .A(n73), .Z(n3597) );
  CNIVXL U5341 ( .A(n73), .Z(n3602) );
  CNIVXL U5342 ( .A(n79), .Z(n3628) );
  CNIVXL U5343 ( .A(n73), .Z(n3595) );
  CNIVXL U5344 ( .A(n79), .Z(n3632) );
  CNIVXL U5345 ( .A(n79), .Z(n3630) );
  CNIVXL U5346 ( .A(n73), .Z(n3598) );
  CNIVXL U5347 ( .A(n73), .Z(n3574) );
  CNIVXL U5348 ( .A(n79), .Z(n3608) );
  CNIVXL U5349 ( .A(n73), .Z(n3600) );
  CNIVXL U5350 ( .A(n73), .Z(n3577) );
  CNIVXL U5351 ( .A(n73), .Z(n3578) );
  CNIVXL U5352 ( .A(n73), .Z(n3599) );
  CNIVXL U5353 ( .A(n73), .Z(n3585) );
  CNIVXL U5354 ( .A(n73), .Z(n3583) );
  CNIVXL U5355 ( .A(n79), .Z(n3626) );
  CNIVXL U5356 ( .A(n73), .Z(n3601) );
  CNIVXL U5357 ( .A(n73), .Z(n3586) );
  CNIVXL U5358 ( .A(n73), .Z(n3596) );
  CNIVXL U5359 ( .A(n73), .Z(n3594) );
  CNIVXL U5360 ( .A(n79), .Z(n3621) );
  CNIVXL U5361 ( .A(n79), .Z(n3611) );
  CNIVXL U5362 ( .A(n79), .Z(n3622) );
  CNIVXL U5363 ( .A(n79), .Z(n3627) );
  CNIVXL U5364 ( .A(n73), .Z(n3575) );
  CNIVXL U5365 ( .A(n73), .Z(n3572) );
  CNIVXL U5366 ( .A(n73), .Z(n3593) );
  CNIVXL U5367 ( .A(n79), .Z(n3607) );
  CNIVXL U5368 ( .A(n79), .Z(n3614) );
  CNIVXL U5369 ( .A(n73), .Z(n3587) );
  CNIVXL U5370 ( .A(n73), .Z(n3588) );
  CNIVXL U5371 ( .A(n73), .Z(n3592) );
  CNIVXL U5372 ( .A(n79), .Z(n3616) );
  CNIVXL U5373 ( .A(n79), .Z(n3623) );
  CNIVXL U5374 ( .A(n79), .Z(n3617) );
  CNIVXL U5375 ( .A(n79), .Z(n3624) );
  CNIVXL U5376 ( .A(n79), .Z(n3625) );
  CNIVXL U5377 ( .A(n79), .Z(n3639) );
  CNIVXL U5378 ( .A(n73), .Z(n3582) );
  CNIVXL U5379 ( .A(n73), .Z(n3581) );
  CNIVXL U5380 ( .A(n73), .Z(n3589) );
  CNIVXL U5381 ( .A(n73), .Z(n3590) );
  CNIVXL U5382 ( .A(n79), .Z(n3615) );
  CNIVXL U5383 ( .A(n73), .Z(n3571) );
  CNIVXL U5384 ( .A(n73), .Z(n3591) );
  CNIVXL U5385 ( .A(n73), .Z(n3580) );
  CNIVXL U5386 ( .A(n73), .Z(n3579) );
  CNIVX2 U5387 ( .A(n75), .Z(n3898) );
  CNR2X1 U5388 ( .A(n4714), .B(n3758), .Z(n4793) );
  CNR2X1 U5389 ( .A(n4734), .B(n3759), .Z(n4803) );
  CNR2XL U5390 ( .A(n5181), .B(n3760), .Z(n5248) );
  CND2IXL U5391 ( .B(n5350), .A(n3737), .Z(n5638) );
  CND2IXL U5392 ( .B(n5913), .A(n3740), .Z(n6143) );
  CNIVX1 U5393 ( .A(n3217), .Z(n3689) );
  CNIVX1 U5394 ( .A(n3217), .Z(n3695) );
  CNIVX1 U5395 ( .A(n3217), .Z(n3683) );
  CNIVX1 U5396 ( .A(n3217), .Z(n3688) );
  CNIVX1 U5397 ( .A(n3217), .Z(n3687) );
  CNIVX1 U5398 ( .A(n3217), .Z(n3690) );
  CNIVX1 U5399 ( .A(n3217), .Z(n3684) );
  CNIVX1 U5400 ( .A(n3217), .Z(n3685) );
  CNIVX1 U5401 ( .A(n3217), .Z(n3693) );
  CNIVX1 U5402 ( .A(n3217), .Z(n3697) );
  CNIVX1 U5403 ( .A(n3217), .Z(n3686) );
  CNIVX1 U5404 ( .A(n3217), .Z(n3696) );
  CNIVX1 U5405 ( .A(n3217), .Z(n3694) );
  CNIVX1 U5406 ( .A(n3217), .Z(n3691) );
  CNIVX1 U5407 ( .A(n3217), .Z(n3698) );
  CNIVX1 U5408 ( .A(n3217), .Z(n3692) );
  CNR2XL U5409 ( .A(n3835), .B(n5212), .Z(N20) );
  CMX2X1 U5410 ( .A0(N7259), .A1(N7258), .S(n3870), .Z(n12693) );
  CMX2XL U5411 ( .A0(N7281), .A1(N7280), .S(n3876), .Z(n12618) );
  CNR2XL U5412 ( .A(n3170), .B(n3221), .Z(n3248) );
  CNR2XL U5413 ( .A(n3170), .B(n3221), .Z(n3249) );
  CNR2XL U5414 ( .A(n3170), .B(n3221), .Z(n74) );
  CND8X1 U5415 ( .A(n3755), .B(n4227), .C(n4437), .D(n3188), .E(n4436), .F(
        n4387), .G(n4400), .H(n3751), .Z(n3170) );
  CMXI2XL U5416 ( .A0(n4624), .A1(n4627), .S(n4214), .Z(n4657) );
  CMXI2X1 U5417 ( .A0(n12169), .A1(n12196), .S(n3452), .Z(N6007) );
  CNR2XL U5418 ( .A(n3509), .B(n12718), .Z(N9301) );
  CNR2XL U5419 ( .A(n3270), .B(n9646), .Z(N6179) );
  CNR2XL U5420 ( .A(n3436), .B(n9645), .Z(N6178) );
  CNR2XL U5421 ( .A(n3439), .B(n12717), .Z(N9300) );
  CNIVX1 U5422 ( .A(n4008), .Z(n4193) );
  CNR2X1 U5423 ( .A(n4706), .B(n3761), .Z(n4789) );
  CNR2XL U5424 ( .A(n4569), .B(n3761), .Z(n6218) );
  CMX2X1 U5425 ( .A0(N7269), .A1(N7268), .S(n3872), .Z(n12667) );
  CMX2X1 U5426 ( .A0(N7285), .A1(N7284), .S(n3864), .Z(n15677) );
  CMX2X1 U5427 ( .A0(N7270), .A1(N7269), .S(n3877), .Z(n12673) );
  CMX2XL U5428 ( .A0(N7259), .A1(N7258), .S(n4287), .Z(n9621) );
  CMX2XL U5429 ( .A0(N7628), .A1(N7627), .S(n3865), .Z(n11466) );
  CNR2X1 U5430 ( .A(n3822), .B(n5425), .Z(n3252) );
  CNR2XL U5431 ( .A(n3815), .B(n4762), .Z(N156) );
  CND2XL U5432 ( .A(n4860), .B(n3728), .Z(n4717) );
  CNR2X1 U5433 ( .A(n5422), .B(n3833), .Z(n3255) );
  CNR2X1 U5434 ( .A(n5415), .B(n3818), .Z(n3258) );
  CNR2X1 U5435 ( .A(n3817), .B(n5423), .Z(n3254) );
  CNR2X1 U5436 ( .A(n3819), .B(n5421), .Z(n3256) );
  CNR2X1 U5437 ( .A(n5414), .B(n3833), .Z(n3259) );
  CNR2X1 U5438 ( .A(n5420), .B(n3820), .Z(n3257) );
  CEOX1 U5439 ( .A(n3265), .B(mem_data1[297]), .Z(N7982) );
  CNR2X1 U5440 ( .A(n3843), .B(n3705), .Z(n3265) );
  CNR2X1 U5441 ( .A(n3839), .B(n3713), .Z(n3264) );
  CMXI2X1 U5442 ( .A0(n4615), .A1(n4614), .S(n4217), .Z(n4671) );
  CNR2IX1 U5443 ( .B(n4655), .A(n3206), .Z(n4827) );
  CNR2IX1 U5444 ( .B(n4758), .A(n3201), .Z(n4821) );
  CMXI2X1 U5445 ( .A0(n12652), .A1(n9638), .S(n3500), .Z(N6164) );
  CMXI2X1 U5446 ( .A0(n12362), .A1(n12389), .S(n3440), .Z(N6064) );
  CMXI2X1 U5447 ( .A0(n12359), .A1(n12386), .S(n3440), .Z(N6063) );
  CMXI2X1 U5448 ( .A0(n12145), .A1(n12169), .S(n3450), .Z(N5999) );
  CMXI2X1 U5449 ( .A0(n12617), .A1(n12643), .S(n3445), .Z(N6143) );
  CMXI2X1 U5450 ( .A0(n12621), .A1(n12645), .S(n3502), .Z(N6144) );
  CMXI2X1 U5451 ( .A0(n11582), .A1(n11609), .S(n3434), .Z(N5831) );
  CMXI2X1 U5452 ( .A0(n11576), .A1(n11600), .S(n3434), .Z(N5829) );
  CMXI2X1 U5453 ( .A0(n11567), .A1(n11594), .S(n3434), .Z(N5827) );
  CMXI2X1 U5454 ( .A0(n11561), .A1(n11588), .S(n3434), .Z(N5825) );
  CMXI2X1 U5455 ( .A0(n11579), .A1(n11606), .S(n3434), .Z(N5830) );
  CMXI2X1 U5456 ( .A0(n11573), .A1(n11597), .S(n3434), .Z(N5828) );
  CMXI2X1 U5457 ( .A0(n11564), .A1(n11591), .S(n3434), .Z(N5826) );
  CMXI2X1 U5458 ( .A0(n11585), .A1(n11612), .S(n3434), .Z(N5832) );
  CMXI2X1 U5459 ( .A0(n11486), .A1(n11513), .S(n3430), .Z(N5802) );
  CMXI2X1 U5460 ( .A0(n11483), .A1(n11510), .S(n3430), .Z(N5801) );
  CMXI2X1 U5461 ( .A0(n11489), .A1(n11516), .S(n3430), .Z(N5803) );
  CND2X1 U5462 ( .A(n5153), .B(n3199), .Z(n5220) );
  CMX2X1 U5463 ( .A0(n5137), .A1(n5207), .S(n3207), .Z(n5266) );
  CMX2X1 U5464 ( .A0(n5134), .A1(n5205), .S(n3203), .Z(n5264) );
  CIVXL U5465 ( .A(n15075), .Z(n4426) );
  CIVXL U5466 ( .A(n14407), .Z(n4427) );
  CND2IXL U5467 ( .B(n12707), .A(n3799), .Z(n12718) );
  CND2IXL U5468 ( .B(n9635), .A(n3218), .Z(n9646) );
  CND2IXL U5469 ( .B(n12705), .A(n3785), .Z(n12717) );
  CND2IXL U5470 ( .B(n9633), .A(n3218), .Z(n9645) );
  CND2IXL U5471 ( .B(n12709), .A(n3801), .Z(n12719) );
  CND2IXL U5472 ( .B(n9637), .A(n3782), .Z(n9647) );
  CND2IXL U5473 ( .B(n12711), .A(n3800), .Z(n12720) );
  CNR2XL U5474 ( .A(n3439), .B(n12716), .Z(N9299) );
  CNR2XL U5475 ( .A(n3270), .B(n12715), .Z(N9298) );
  CNR2XL U5476 ( .A(n3270), .B(n12714), .Z(N9297) );
  CNR2XL U5477 ( .A(n3270), .B(n12713), .Z(N9296) );
  CMX2XL U5478 ( .A0(n5248), .A1(n5182), .S(n3200), .Z(n5286) );
  CMX2XL U5479 ( .A0(n5143), .A1(n5213), .S(n3215), .Z(n5268) );
  COR2XL U5480 ( .A(n3604), .B(n3682), .Z(n3250) );
  CNIVXL U5481 ( .A(n4008), .Z(n4198) );
  CMXI2X1 U5482 ( .A0(n4650), .A1(n4649), .S(n4226), .Z(n4728) );
  CNR2X1 U5483 ( .A(n4747), .B(n3765), .Z(n4811) );
  CNR2X1 U5484 ( .A(n5175), .B(n3761), .Z(n5242) );
  CNR2X1 U5485 ( .A(n4689), .B(n3762), .Z(n4751) );
  CNR2X1 U5486 ( .A(n4701), .B(n3762), .Z(n4757) );
  CNR2X1 U5487 ( .A(n6172), .B(n3758), .Z(n6206) );
  CND2X1 U5488 ( .A(n5290), .B(n3738), .Z(n5463) );
  CND2X1 U5489 ( .A(n4882), .B(n3738), .Z(n6019) );
  CND2X1 U5490 ( .A(n5708), .B(n4221), .Z(n5745) );
  CND2X1 U5491 ( .A(n4659), .B(n3894), .Z(n4697) );
  CND2X1 U5492 ( .A(n4951), .B(n3892), .Z(n5003) );
  CND2X1 U5493 ( .A(n4817), .B(n3740), .Z(n4926) );
  CND2IX1 U5494 ( .B(n5208), .A(n3726), .Z(n5311) );
  CNR2XL U5495 ( .A(n4726), .B(n3761), .Z(n4799) );
  CNR2XL U5496 ( .A(n4710), .B(n3759), .Z(n4791) );
  CNR2XL U5497 ( .A(n4730), .B(n3758), .Z(n4801) );
  CMXI2X1 U5498 ( .A0(n13740), .A1(n13739), .S(n4178), .Z(n13741) );
  CND2XL U5499 ( .A(n5102), .B(n3190), .Z(n5121) );
  CND2IXL U5500 ( .B(n5194), .A(n3730), .Z(n5296) );
  CND2IXL U5501 ( .B(n5354), .A(n3737), .Z(n5653) );
  CND2IXL U5502 ( .B(n5917), .A(n3739), .Z(n6149) );
  CND2IXL U5503 ( .B(n5907), .A(n3731), .Z(n6134) );
  CND2IXL U5504 ( .B(n5909), .A(n3731), .Z(n6137) );
  CND2IXL U5505 ( .B(n6238), .A(n3726), .Z(n6340) );
  CND2IXL U5506 ( .B(n6240), .A(n3727), .Z(n6342) );
  CND2IXL U5507 ( .B(n5757), .A(n3728), .Z(n5860) );
  CND2IXL U5508 ( .B(n5903), .A(n3732), .Z(n6128) );
  CND2IXL U5509 ( .B(n5905), .A(n3740), .Z(n6131) );
  CND2IXL U5510 ( .B(n5352), .A(n3732), .Z(n5646) );
  CND2IXL U5511 ( .B(n5348), .A(n3736), .Z(n5631) );
  CND2XL U5512 ( .A(n9630), .B(n4010), .Z(n9639) );
  CANR2XL U5513 ( .A(N3105), .B(n3592), .C(n3200), .D(n3637), .Z(n2114) );
  CND2X1 U5514 ( .A(n4400), .B(n5604), .Z(n4543) );
  CNR2XL U5515 ( .A(n4920), .B(n4220), .Z(n4939) );
  CMX2X1 U5516 ( .A0(N7273), .A1(N7272), .S(n3878), .Z(n12665) );
  CND2XL U5517 ( .A(n4589), .B(n3194), .Z(n4633) );
  CND2XL U5518 ( .A(n4475), .B(n3190), .Z(n4501) );
  CND2XL U5519 ( .A(n5671), .B(n3192), .Z(n5688) );
  CND2XL U5520 ( .A(n5107), .B(n3188), .Z(n5125) );
  CND2XL U5521 ( .A(n4935), .B(n4407), .Z(n6062) );
  CND2XL U5522 ( .A(n6041), .B(n4410), .Z(n6047) );
  CND2XL U5523 ( .A(n6037), .B(n4413), .Z(n6042) );
  CND2XL U5524 ( .A(n6032), .B(n4413), .Z(n6038) );
  CND2XL U5525 ( .A(n5604), .B(n4411), .Z(n5612) );
  CAN2XL U5526 ( .A(N7256), .B(n3886), .Z(n12702) );
  CMX2XL U5527 ( .A0(N7261), .A1(N7260), .S(n4287), .Z(n9615) );
  CMX2XL U5528 ( .A0(N7261), .A1(N7260), .S(n3868), .Z(n12687) );
  CMX2XL U5529 ( .A0(N7264), .A1(N7263), .S(n4287), .Z(n9604) );
  CMX2XL U5530 ( .A0(N7265), .A1(N7264), .S(n3881), .Z(n12669) );
  CMX2XL U5531 ( .A0(N7265), .A1(N7264), .S(n4288), .Z(n9597) );
  CMX2XL U5532 ( .A0(N7260), .A1(N7259), .S(n4287), .Z(n9619) );
  CMX2XL U5533 ( .A0(N7269), .A1(N7268), .S(n4288), .Z(n9595) );
  CMX2XL U5534 ( .A0(N7285), .A1(N7284), .S(n3872), .Z(n12606) );
  CMX2XL U5535 ( .A0(N7268), .A1(N7267), .S(n4287), .Z(n9602) );
  CMX2XL U5536 ( .A0(N7284), .A1(N7283), .S(n3873), .Z(n12609) );
  CMX2XL U5537 ( .A0(N7270), .A1(N7269), .S(n4287), .Z(n9601) );
  CMX2XL U5538 ( .A0(N7286), .A1(N7285), .S(n3871), .Z(n12603) );
  CMX2XL U5539 ( .A0(N7282), .A1(N7281), .S(n3875), .Z(n12615) );
  CMX2XL U5540 ( .A0(N7262), .A1(N7261), .S(n3872), .Z(n12683) );
  CMX2XL U5541 ( .A0(N7262), .A1(N7261), .S(n4287), .Z(n9611) );
  CMX2XL U5542 ( .A0(N7263), .A1(N7262), .S(n4287), .Z(n9607) );
  CMX2XL U5543 ( .A0(N7267), .A1(N7266), .S(n4288), .Z(n9596) );
  CMX2XL U5544 ( .A0(N7266), .A1(N7265), .S(n3878), .Z(n12675) );
  CMX2XL U5545 ( .A0(N7266), .A1(N7265), .S(n4287), .Z(n9603) );
  CMX2XL U5546 ( .A0(N7287), .A1(N7286), .S(n3877), .Z(n12600) );
  CMX2XL U5547 ( .A0(N7283), .A1(N7282), .S(n3874), .Z(n12612) );
  CMX2XL U5548 ( .A0(N7271), .A1(N7270), .S(n4288), .Z(n9594) );
  CMX2XL U5549 ( .A0(N7258), .A1(N7257), .S(n4285), .Z(n9624) );
  CMX2XL U5550 ( .A0(N7257), .A1(N7256), .S(n4286), .Z(n9627) );
  CMX2XL U5551 ( .A0(N7257), .A1(N7256), .S(n3864), .Z(n12699) );
  CANR2XL U5552 ( .A(N2428), .B(n3582), .C(n3617), .D(N7927), .Z(n1048) );
  CIVX2 U5553 ( .A(lenin0[1]), .Z(n4428) );
  CNR2X1 U5554 ( .A(n3852), .B(n5986), .Z(N24) );
  CNR2XL U5555 ( .A(n3837), .B(n4881), .Z(N19) );
  CNR2X1 U5556 ( .A(n3817), .B(n4784), .Z(N160) );
  CND2XL U5557 ( .A(n4822), .B(n3726), .Z(n4611) );
  CND2XL U5558 ( .A(n4835), .B(n3722), .Z(n4661) );
  CAN2XL U5559 ( .A(datain0[27]), .B(n4389), .Z(n5625) );
  CAN2XL U5560 ( .A(datain0[23]), .B(n4389), .Z(n5597) );
  CAN2XL U5561 ( .A(datain0[22]), .B(n4389), .Z(n5590) );
  CAN2XL U5562 ( .A(datain0[21]), .B(n4389), .Z(n5583) );
  CAN2XL U5563 ( .A(datain0[20]), .B(n4389), .Z(n5576) );
  CND2XL U5564 ( .A(n2112), .B(n2113), .Z(N10354) );
  CND2X1 U5565 ( .A(n5120), .B(n3205), .Z(n5198) );
  CMXI2XL U5566 ( .A0(n4622), .A1(n4625), .S(n4212), .Z(n4658) );
  CMXI2XL U5567 ( .A0(n4625), .A1(n4624), .S(n4219), .Z(n4677) );
  CND2X1 U5568 ( .A(n5124), .B(n3207), .Z(n5200) );
  CMXI2XL U5569 ( .A0(n12389), .A1(n12416), .S(n3439), .Z(N6072) );
  CNR2IXL U5570 ( .B(n4800), .A(n3202), .Z(n4866) );
  CNR2IXL U5571 ( .B(n4765), .A(n3200), .Z(n4833) );
  CNR2IXL U5572 ( .B(n4761), .A(n3212), .Z(n4824) );
  CNR2IXL U5573 ( .B(n4705), .A(n3210), .Z(n4829) );
  CND2XL U5574 ( .A(n5788), .B(n3202), .Z(n5890) );
  CND2XL U5575 ( .A(n5792), .B(n3204), .Z(n5894) );
  CMX2XL U5576 ( .A0(n5146), .A1(n5215), .S(n3209), .Z(n5269) );
  CAN2XL U5577 ( .A(n5187), .B(n3206), .Z(n5290) );
  CANR2XL U5578 ( .A(N6226), .B(n2105), .C(n3759), .D(n3898), .Z(n2117) );
  CND2XL U5579 ( .A(n2116), .B(n2117), .Z(N10352) );
  CANR2XL U5580 ( .A(N3108), .B(n3592), .C(N2074), .D(n3637), .Z(n2108) );
  CANR2XL U5581 ( .A(N6228), .B(n2105), .C(n3898), .D(n3726), .Z(n2113) );
  CANR2XL U5582 ( .A(N6229), .B(n2105), .C(n3898), .D(n3818), .Z(n2111) );
  CANR2XL U5583 ( .A(N3107), .B(n3592), .C(N2073), .D(n3637), .Z(n2110) );
  CND2XL U5584 ( .A(n2118), .B(n2119), .Z(N10351) );
  CANR2XL U5585 ( .A(N6225), .B(n2105), .C(n3891), .D(n3898), .Z(n2119) );
  CIVX1 U5586 ( .A(n3569), .Z(n3533) );
  CNIVXL U5587 ( .A(n4437), .Z(n4216) );
  CNIVXL U5588 ( .A(n4437), .Z(n4220) );
  CNIVXL U5589 ( .A(n4437), .Z(n4213) );
  CNIVXL U5590 ( .A(n4437), .Z(n4212) );
  CMXI2XL U5591 ( .A0(n5102), .A1(n5092), .S(n3190), .Z(n5113) );
  CMXI2XL U5592 ( .A0(n4677), .A1(n4680), .S(n4221), .Z(n4716) );
  CMXI2XL U5593 ( .A0(n4656), .A1(n4658), .S(n4223), .Z(n4696) );
  CMXI2XL U5594 ( .A0(n13403), .A1(n13402), .S(n4185), .Z(n13404) );
  CNR2XL U5595 ( .A(n3763), .B(n5074), .Z(n5146) );
  CNR2XL U5596 ( .A(n5031), .B(n3762), .Z(n5128) );
  CNR2XL U5597 ( .A(n5010), .B(n3763), .Z(n5116) );
  CNR2XL U5598 ( .A(n4996), .B(n3764), .Z(n5106) );
  CNR2XL U5599 ( .A(n4700), .B(n3760), .Z(n4787) );
  CNR2XL U5600 ( .A(n4533), .B(n3761), .Z(n6212) );
  CNR2XL U5601 ( .A(n3764), .B(n5067), .Z(n5143) );
  CND2XL U5602 ( .A(n3721), .B(n4876), .Z(n5568) );
  CND2XL U5603 ( .A(n4883), .B(n3731), .Z(n6036) );
  CND2XL U5604 ( .A(n4884), .B(n3734), .Z(n6085) );
  CND2XL U5605 ( .A(n5699), .B(n4221), .Z(n5738) );
  CND2XL U5606 ( .A(n5705), .B(n4221), .Z(n5743) );
  CND2XL U5607 ( .A(n5141), .B(n4222), .Z(n5179) );
  CND2XL U5608 ( .A(n4642), .B(n4223), .Z(n4722) );
  CND2XL U5609 ( .A(n4813), .B(n3739), .Z(n4917) );
  CND2XL U5610 ( .A(n4821), .B(n3739), .Z(n4934) );
  CND2IXL U5611 ( .B(n5865), .A(n3732), .Z(n6050) );
  CND2IXL U5612 ( .B(n5878), .A(n3740), .Z(n6080) );
  CND2IXL U5613 ( .B(n5873), .A(n3739), .Z(n6071) );
  CND2IXL U5614 ( .B(n5789), .A(n3725), .Z(n5891) );
  CND2IXL U5615 ( .B(n5901), .A(n3733), .Z(n6124) );
  CND2IXL U5616 ( .B(n5899), .A(n3734), .Z(n6120) );
  CND2IXL U5617 ( .B(n5896), .A(n3738), .Z(n6116) );
  CND2IXL U5618 ( .B(n5892), .A(n3735), .Z(n6108) );
  CND2IXL U5619 ( .B(n5888), .A(n3734), .Z(n6100) );
  CND2IXL U5620 ( .B(n5886), .A(n3734), .Z(n6096) );
  CND2IXL U5621 ( .B(n5778), .A(n3725), .Z(n5881) );
  CND2IXL U5622 ( .B(n5776), .A(n3727), .Z(n5879) );
  CND2IXL U5623 ( .B(n5774), .A(n3725), .Z(n5876) );
  CND2IXL U5624 ( .B(n5345), .A(n3737), .Z(n5624) );
  CND2IXL U5625 ( .B(n5780), .A(n3726), .Z(n5883) );
  CND2IXL U5626 ( .B(n5772), .A(n3727), .Z(n5874) );
  CND2IXL U5627 ( .B(n5770), .A(n3728), .Z(n5872) );
  CND2IXL U5628 ( .B(n5766), .A(n3722), .Z(n5868) );
  CND2IXL U5629 ( .B(n5764), .A(n3724), .Z(n5866) );
  CND2IXL U5630 ( .B(n5761), .A(n3730), .Z(n5864) );
  CND2IXL U5631 ( .B(n5343), .A(n3740), .Z(n5617) );
  CND2IXL U5632 ( .B(n5341), .A(n3735), .Z(n5610) );
  CND2IXL U5633 ( .B(n5206), .A(n3726), .Z(n5309) );
  CND2IXL U5634 ( .B(n5200), .A(n3727), .Z(n5302) );
  CANR2XL U5635 ( .A(N6231), .B(n2105), .C(n3898), .D(n4400), .Z(n2107) );
  CND2XL U5636 ( .A(n2106), .B(n2107), .Z(N10357) );
  CND2XL U5637 ( .A(n2114), .B(n2115), .Z(N10353) );
  CND2XL U5638 ( .A(n2120), .B(n2121), .Z(N10350) );
  CANR2XL U5639 ( .A(N6224), .B(n2105), .C(n3896), .D(n3898), .Z(n2121) );
  CNIVXL U5640 ( .A(n3249), .Z(n3677) );
  CNIVXL U5641 ( .A(n3248), .Z(n3674) );
  CNIVXL U5642 ( .A(n3249), .Z(n3665) );
  CNIVXL U5643 ( .A(n3248), .Z(n3641) );
  CNIVXL U5644 ( .A(n3249), .Z(n3642) );
  CNIVXL U5645 ( .A(n3248), .Z(n3643) );
  CNIVXL U5646 ( .A(n3249), .Z(n3644) );
  CNIVXL U5647 ( .A(n3249), .Z(n3682) );
  CNIVXL U5648 ( .A(n3756), .Z(n3761) );
  CNIVXL U5649 ( .A(n3756), .Z(n3758) );
  CND2XL U5650 ( .A(\r347/carry [8]), .B(n4389), .Z(n3267) );
  CNR2XL U5651 ( .A(n4613), .B(n3896), .Z(n4648) );
  CMX2XL U5652 ( .A0(N7527), .A1(N7526), .S(n3872), .Z(n11806) );
  CMX2XL U5653 ( .A0(N7280), .A1(N7279), .S(n3881), .Z(n15693) );
  CMX2XL U5654 ( .A0(N7272), .A1(N7271), .S(n3863), .Z(n12672) );
  CMX2XL U5655 ( .A0(N7279), .A1(N7278), .S(n4288), .Z(n12619) );
  CMX2XL U5656 ( .A0(N7280), .A1(N7279), .S(n3877), .Z(n12622) );
  CMX2XL U5657 ( .A0(N7273), .A1(N7272), .S(n4288), .Z(n9593) );
  CMX2XL U5658 ( .A0(N7756), .A1(N7755), .S(n4250), .Z(n11042) );
  CMX2XL U5659 ( .A0(N7272), .A1(N7271), .S(n4287), .Z(n9600) );
  CMX2XL U5660 ( .A0(N7564), .A1(N7563), .S(n3864), .Z(n11683) );
  CMX2XL U5661 ( .A0(N7692), .A1(N7691), .S(n3870), .Z(n11252) );
  CNIVXL U5662 ( .A(n3756), .Z(n3760) );
  CNIVXL U5663 ( .A(n3756), .Z(n3759) );
  CNIVXL U5664 ( .A(n3249), .Z(n3671) );
  CNIVXL U5665 ( .A(n3248), .Z(n3673) );
  CNIVXL U5666 ( .A(n3248), .Z(n3672) );
  CNIVXL U5667 ( .A(n3249), .Z(n3663) );
  CNIVXL U5668 ( .A(n3249), .Z(n3661) );
  CNIVXL U5669 ( .A(n3249), .Z(n3660) );
  CNIVXL U5670 ( .A(n3248), .Z(n3662) );
  CNIVXL U5671 ( .A(n3248), .Z(n3669) );
  CNIVXL U5672 ( .A(n3249), .Z(n3668) );
  CNIVXL U5673 ( .A(n3248), .Z(n3670) );
  CNIVXL U5674 ( .A(n3249), .Z(n3667) );
  CNIVXL U5675 ( .A(n3248), .Z(n3664) );
  CNIVXL U5676 ( .A(n3249), .Z(n3666) );
  CNIVXL U5677 ( .A(n3248), .Z(n3652) );
  CNIVXL U5678 ( .A(n3249), .Z(n3653) );
  CNIVXL U5679 ( .A(n3248), .Z(n3654) );
  CNIVXL U5680 ( .A(n3249), .Z(n3655) );
  CNIVXL U5681 ( .A(n3248), .Z(n3656) );
  CNIVXL U5682 ( .A(n3249), .Z(n3657) );
  CNIVXL U5683 ( .A(n3248), .Z(n3658) );
  CNIVXL U5684 ( .A(n3248), .Z(n3659) );
  CND2XL U5685 ( .A(n2122), .B(n2123), .Z(N10349) );
  CANR2XL U5686 ( .A(mem_data1[1020]), .B(n3898), .C(N9300), .D(n3674), .Z(
        n2135) );
  CANR2XL U5687 ( .A(mem_data1[1019]), .B(n3898), .C(N9299), .D(n3674), .Z(
        n2138) );
  CANR2XL U5688 ( .A(mem_data1[1018]), .B(n3898), .C(N9298), .D(n3674), .Z(
        n2141) );
  CANR2XL U5689 ( .A(mem_data1[1017]), .B(n3898), .C(N9297), .D(n3674), .Z(
        n2144) );
  CANR2XL U5690 ( .A(mem_data1[1016]), .B(n3898), .C(N9296), .D(n3674), .Z(
        n2147) );
  CANR2XL U5691 ( .A(mem_data1[1015]), .B(n3898), .C(N9295), .D(n3674), .Z(
        n2150) );
  CANR2XL U5692 ( .A(mem_data1[1014]), .B(n3898), .C(N9294), .D(n3674), .Z(
        n2153) );
  CANR2XL U5693 ( .A(mem_data1[1013]), .B(n3898), .C(N9293), .D(n3674), .Z(
        n2156) );
  CANR2XL U5694 ( .A(mem_data1[1011]), .B(n3898), .C(N9291), .D(n3675), .Z(
        n2162) );
  CANR2XL U5695 ( .A(mem_data1[1010]), .B(n3898), .C(N9290), .D(n3675), .Z(
        n2165) );
  CANR2XL U5696 ( .A(mem_data1[1009]), .B(n3898), .C(N9289), .D(n3675), .Z(
        n2168) );
  CANR2XL U5697 ( .A(mem_data1[1008]), .B(n3898), .C(N9288), .D(n3675), .Z(
        n2171) );
  CANR2XL U5698 ( .A(N3083), .B(n3593), .C(n3627), .D(N7272), .Z(n2176) );
  CANR2XL U5699 ( .A(mem_data1[1007]), .B(n3898), .C(N9287), .D(n3675), .Z(
        n2174) );
  CANR2XL U5700 ( .A(N3082), .B(n3593), .C(n3627), .D(N7273), .Z(n2179) );
  CND2XL U5701 ( .A(N6164), .B(n3691), .Z(n2178) );
  CANR2XL U5702 ( .A(mem_data1[1006]), .B(n3898), .C(N9286), .D(n3675), .Z(
        n2177) );
  CANR2XL U5703 ( .A(mem_data1[1022]), .B(n3898), .C(N9302), .D(n3674), .Z(
        n2129) );
  CANR2XL U5704 ( .A(mem_data1[1023]), .B(n3898), .C(N9303), .D(n3674), .Z(
        n2126) );
  CND2XL U5705 ( .A(N5450), .B(n3691), .Z(n1227) );
  CANR2XL U5706 ( .A(mem_data1[292]), .B(n3898), .C(N8572), .D(n3679), .Z(
        n1226) );
  CND2XL U5707 ( .A(N5451), .B(n3688), .Z(n1224) );
  CANR2XL U5708 ( .A(mem_data1[293]), .B(n3898), .C(N8573), .D(n3679), .Z(
        n1223) );
  CND2XL U5709 ( .A(N5461), .B(n3686), .Z(n1194) );
  CANR2XL U5710 ( .A(mem_data1[303]), .B(n3898), .C(N8583), .D(n3679), .Z(
        n1193) );
  CND2XL U5711 ( .A(N5463), .B(n3693), .Z(n1188) );
  CANR2XL U5712 ( .A(mem_data1[305]), .B(n3898), .C(N8585), .D(n3679), .Z(
        n1187) );
  CND2XL U5713 ( .A(N5574), .B(n3689), .Z(n855) );
  CANR2XL U5714 ( .A(N2492), .B(n3580), .C(n3616), .D(N7863), .Z(n856) );
  CND2XL U5715 ( .A(N5448), .B(n3688), .Z(n1233) );
  CANR2XL U5716 ( .A(mem_data1[290]), .B(n3898), .C(N8570), .D(n3679), .Z(
        n1232) );
  CND2XL U5717 ( .A(N5404), .B(n3688), .Z(n1365) );
  CANR2XL U5718 ( .A(mem_data1[246]), .B(n3898), .C(N8526), .D(n3680), .Z(
        n1364) );
  CND2XL U5719 ( .A(N5603), .B(n3687), .Z(n768) );
  CANR2XL U5720 ( .A(mem_data1[445]), .B(n3898), .C(N8725), .D(n3679), .Z(n767) );
  CND2XL U5721 ( .A(N5649), .B(n3686), .Z(n630) );
  CANR2XL U5722 ( .A(mem_data1[491]), .B(n3898), .C(N8771), .D(n3681), .Z(n629) );
  CND2XL U5723 ( .A(N5651), .B(n3686), .Z(n624) );
  CANR2XL U5724 ( .A(N2569), .B(n3570), .C(n3606), .D(N7786), .Z(n625) );
  CND2XL U5725 ( .A(N5650), .B(n3686), .Z(n627) );
  CANR2XL U5726 ( .A(mem_data1[492]), .B(n3898), .C(N8772), .D(n3681), .Z(n626) );
  CND2XL U5727 ( .A(N5473), .B(n3696), .Z(n1158) );
  CANR2XL U5728 ( .A(mem_data1[315]), .B(n3898), .C(N8595), .D(n3680), .Z(
        n1157) );
  CND2XL U5729 ( .A(N5475), .B(n3698), .Z(n1152) );
  CANR2XL U5730 ( .A(mem_data1[317]), .B(n3898), .C(N8597), .D(n3680), .Z(
        n1151) );
  CND2XL U5731 ( .A(N5590), .B(n3686), .Z(n807) );
  CANR2XL U5732 ( .A(N2508), .B(n3571), .C(n3608), .D(N7847), .Z(n808) );
  CND2XL U5733 ( .A(N5571), .B(n3689), .Z(n864) );
  CANR2XL U5734 ( .A(mem_data1[413]), .B(n3898), .C(N8693), .D(n3681), .Z(n863) );
  CND2XL U5735 ( .A(N5539), .B(n3696), .Z(n960) );
  CANR2XL U5736 ( .A(mem_data1[381]), .B(n3898), .C(N8661), .D(n3681), .Z(n959) );
  CND2XL U5737 ( .A(N5538), .B(n3693), .Z(n963) );
  CANR2XL U5738 ( .A(mem_data1[380]), .B(n3898), .C(N8660), .D(n3681), .Z(n962) );
  CND2XL U5739 ( .A(N5505), .B(n3690), .Z(n1062) );
  CANR2XL U5740 ( .A(N2423), .B(n3582), .C(n3617), .D(N7932), .Z(n1063) );
  CND2XL U5741 ( .A(N5510), .B(n3698), .Z(n1047) );
  CND2XL U5742 ( .A(N5516), .B(n3698), .Z(n1029) );
  CANR2XL U5743 ( .A(mem_data1[358]), .B(n3898), .C(N8638), .D(n3680), .Z(
        n1028) );
  CND2XL U5744 ( .A(N5515), .B(n3689), .Z(n1032) );
  CANR2XL U5745 ( .A(mem_data1[357]), .B(n3898), .C(N8637), .D(n3681), .Z(
        n1031) );
  CND2XL U5746 ( .A(N5537), .B(n3688), .Z(n966) );
  CANR2XL U5747 ( .A(mem_data1[379]), .B(n3898), .C(N8659), .D(n3681), .Z(n965) );
  CANR2XL U5748 ( .A(N3081), .B(n3593), .C(n3627), .D(N7274), .Z(n2182) );
  CND2XL U5749 ( .A(N6163), .B(n3691), .Z(n2181) );
  CANR2XL U5750 ( .A(mem_data1[1005]), .B(n3898), .C(N9285), .D(n3675), .Z(
        n2180) );
  CANR2XL U5751 ( .A(N3080), .B(n3593), .C(n3627), .D(N7275), .Z(n2185) );
  CND2XL U5752 ( .A(N6162), .B(n3685), .Z(n2184) );
  CANR2XL U5753 ( .A(mem_data1[1004]), .B(n3898), .C(N9284), .D(n3675), .Z(
        n2183) );
  CANR2XL U5754 ( .A(N3065), .B(n3595), .C(n3629), .D(N7290), .Z(n2230) );
  CND2XL U5755 ( .A(N6147), .B(n3693), .Z(n2229) );
  CANR2XL U5756 ( .A(mem_data1[989]), .B(n3898), .C(N9269), .D(n3674), .Z(
        n2228) );
  CANR2XL U5757 ( .A(N3064), .B(n3594), .C(n3628), .D(N7291), .Z(n2233) );
  CND2XL U5758 ( .A(N6146), .B(n3693), .Z(n2232) );
  CANR2XL U5759 ( .A(mem_data1[988]), .B(n3898), .C(N9268), .D(n3674), .Z(
        n2231) );
  CANR2XL U5760 ( .A(N3063), .B(n3594), .C(n3628), .D(N7292), .Z(n2236) );
  CND2XL U5761 ( .A(N6145), .B(n3693), .Z(n2235) );
  CANR2XL U5762 ( .A(mem_data1[987]), .B(n3898), .C(N9267), .D(n3674), .Z(
        n2234) );
  CANR2XL U5763 ( .A(N3062), .B(n3594), .C(n3628), .D(N7293), .Z(n2239) );
  CND2XL U5764 ( .A(N6144), .B(n3693), .Z(n2238) );
  CANR2XL U5765 ( .A(mem_data1[986]), .B(n3898), .C(N9266), .D(n3674), .Z(
        n2237) );
  CANR2XL U5766 ( .A(N3061), .B(n3594), .C(n3628), .D(N7294), .Z(n2242) );
  CND2XL U5767 ( .A(N6143), .B(n3693), .Z(n2241) );
  CANR2XL U5768 ( .A(mem_data1[985]), .B(n3898), .C(N9265), .D(n3674), .Z(
        n2240) );
  CANR2XL U5769 ( .A(N3060), .B(n3594), .C(n3628), .D(N7295), .Z(n2245) );
  CANR2XL U5770 ( .A(mem_data1[984]), .B(n3898), .C(N9264), .D(n3674), .Z(
        n2243) );
  CANR2XL U5771 ( .A(N3059), .B(n3594), .C(n3628), .D(N7296), .Z(n2248) );
  CANR2XL U5772 ( .A(mem_data1[983]), .B(n3898), .C(N9263), .D(n3674), .Z(
        n2246) );
  CANR2XL U5773 ( .A(N3058), .B(n3594), .C(n3630), .D(N7297), .Z(n2251) );
  CANR2XL U5774 ( .A(mem_data1[982]), .B(n3898), .C(N9262), .D(n3674), .Z(
        n2249) );
  CND2XL U5775 ( .A(N6115), .B(n3692), .Z(n2325) );
  CANR2XL U5776 ( .A(N3033), .B(n3595), .C(n3629), .D(N7322), .Z(n2326) );
  CANR2XL U5777 ( .A(N3005), .B(n3600), .C(n3634), .D(N7350), .Z(n2410) );
  CND2XL U5778 ( .A(N6087), .B(n3698), .Z(n2409) );
  CANR2XL U5779 ( .A(mem_data1[929]), .B(n3898), .C(N9209), .D(n3674), .Z(
        n2408) );
  CANR2XL U5780 ( .A(N2990), .B(n3600), .C(n3633), .D(N7365), .Z(n2455) );
  CND2XL U5781 ( .A(N6072), .B(n3687), .Z(n2454) );
  CANR2XL U5782 ( .A(mem_data1[914]), .B(n3898), .C(N9194), .D(n3676), .Z(
        n2453) );
  CANR2XL U5783 ( .A(N2989), .B(n3600), .C(n3633), .D(N7366), .Z(n2458) );
  CANR2XL U5784 ( .A(mem_data1[913]), .B(n3898), .C(N9193), .D(n3676), .Z(
        n2456) );
  CANR2XL U5785 ( .A(mem_data1[912]), .B(n3898), .C(N9192), .D(n3676), .Z(
        n2459) );
  CANR2XL U5786 ( .A(N2987), .B(n3599), .C(n3633), .D(N7368), .Z(n2464) );
  CANR2XL U5787 ( .A(mem_data1[911]), .B(n3898), .C(N9191), .D(n3676), .Z(
        n2462) );
  CANR2XL U5788 ( .A(N2986), .B(n3601), .C(n3633), .D(N7369), .Z(n2467) );
  CANR2XL U5789 ( .A(mem_data1[910]), .B(n3898), .C(N9190), .D(n3676), .Z(
        n2465) );
  CANR2XL U5790 ( .A(N2985), .B(n3601), .C(n3633), .D(N7370), .Z(n2470) );
  CANR2XL U5791 ( .A(mem_data1[909]), .B(n3898), .C(N9189), .D(n3676), .Z(
        n2468) );
  CANR2XL U5792 ( .A(N2984), .B(n3601), .C(n3633), .D(N7371), .Z(n2473) );
  CANR2XL U5793 ( .A(mem_data1[908]), .B(n3898), .C(N9188), .D(n3676), .Z(
        n2471) );
  CANR2XL U5794 ( .A(N2983), .B(n3601), .C(n3633), .D(N7372), .Z(n2476) );
  CANR2XL U5795 ( .A(mem_data1[907]), .B(n3898), .C(N9187), .D(n3675), .Z(
        n2474) );
  CANR2XL U5796 ( .A(N2982), .B(n3601), .C(n3610), .D(N7373), .Z(n2479) );
  CND2XL U5797 ( .A(N6064), .B(n3698), .Z(n2478) );
  CANR2XL U5798 ( .A(mem_data1[906]), .B(n3898), .C(N9186), .D(n3675), .Z(
        n2477) );
  CANR2XL U5799 ( .A(N2981), .B(n3601), .C(n3612), .D(N7374), .Z(n2482) );
  CND2XL U5800 ( .A(N6063), .B(n3686), .Z(n2481) );
  CANR2XL U5801 ( .A(mem_data1[905]), .B(n3898), .C(N9185), .D(n3675), .Z(
        n2480) );
  CANR2XL U5802 ( .A(N2980), .B(n3601), .C(n3614), .D(N7375), .Z(n2485) );
  CND2XL U5803 ( .A(N6062), .B(n3694), .Z(n2484) );
  CANR2XL U5804 ( .A(mem_data1[904]), .B(n3898), .C(N9184), .D(n3675), .Z(
        n2483) );
  CANR2XL U5805 ( .A(N2979), .B(n3601), .C(n3631), .D(N7376), .Z(n2488) );
  CND2XL U5806 ( .A(N6061), .B(n3691), .Z(n2487) );
  CANR2XL U5807 ( .A(mem_data1[903]), .B(n3898), .C(N9183), .D(n3675), .Z(
        n2486) );
  CANR2XL U5808 ( .A(N2949), .B(n3574), .C(n3610), .D(N7406), .Z(n2578) );
  CND2XL U5809 ( .A(N6031), .B(n3687), .Z(n2577) );
  CANR2XL U5810 ( .A(mem_data1[873]), .B(n3898), .C(N9153), .D(n3677), .Z(
        n2576) );
  CANR2XL U5811 ( .A(N2948), .B(n3574), .C(n3610), .D(N7407), .Z(n2581) );
  CND2XL U5812 ( .A(N6030), .B(n3688), .Z(n2580) );
  CANR2XL U5813 ( .A(mem_data1[872]), .B(n3898), .C(N9152), .D(n3676), .Z(
        n2579) );
  CANR2XL U5814 ( .A(N2925), .B(n3575), .C(n3612), .D(N7430), .Z(n2650) );
  CND2XL U5815 ( .A(N6007), .B(n3695), .Z(n2649) );
  CANR2XL U5816 ( .A(mem_data1[849]), .B(n3898), .C(N9129), .D(n3661), .Z(
        n2648) );
  CND2XL U5817 ( .A(N6006), .B(n3695), .Z(n2652) );
  CANR2XL U5818 ( .A(mem_data1[848]), .B(n3898), .C(N9128), .D(n3661), .Z(
        n2651) );
  CANR2XL U5819 ( .A(N2923), .B(n3575), .C(n3611), .D(N7432), .Z(n2656) );
  CND2XL U5820 ( .A(N6005), .B(n3695), .Z(n2655) );
  CANR2XL U5821 ( .A(mem_data1[847]), .B(n3898), .C(N9127), .D(n3661), .Z(
        n2654) );
  CANR2XL U5822 ( .A(N2922), .B(n3575), .C(n3611), .D(N7433), .Z(n2659) );
  CND2XL U5823 ( .A(N6004), .B(n3695), .Z(n2658) );
  CANR2XL U5824 ( .A(mem_data1[846]), .B(n3898), .C(N9126), .D(n3662), .Z(
        n2657) );
  CANR2XL U5825 ( .A(N2921), .B(n3575), .C(n3611), .D(N7434), .Z(n2662) );
  CND2XL U5826 ( .A(N6003), .B(n3695), .Z(n2661) );
  CANR2XL U5827 ( .A(mem_data1[845]), .B(n3898), .C(N9125), .D(n3662), .Z(
        n2660) );
  CANR2XL U5828 ( .A(N2920), .B(n3575), .C(n3611), .D(N7435), .Z(n2665) );
  CND2XL U5829 ( .A(N6002), .B(n3694), .Z(n2664) );
  CANR2XL U5830 ( .A(mem_data1[844]), .B(n3898), .C(N9124), .D(n3662), .Z(
        n2663) );
  CANR2XL U5831 ( .A(N2919), .B(n3575), .C(n3611), .D(N7436), .Z(n2668) );
  CND2XL U5832 ( .A(N6001), .B(n3696), .Z(n2667) );
  CANR2XL U5833 ( .A(mem_data1[843]), .B(n3898), .C(N9123), .D(n3662), .Z(
        n2666) );
  CANR2XL U5834 ( .A(N2918), .B(n3575), .C(n3611), .D(N7437), .Z(n2671) );
  CND2XL U5835 ( .A(N6000), .B(n3695), .Z(n2670) );
  CANR2XL U5836 ( .A(mem_data1[842]), .B(n3898), .C(N9122), .D(n3662), .Z(
        n2669) );
  CANR2XL U5837 ( .A(N2917), .B(n3575), .C(n3611), .D(N7438), .Z(n2674) );
  CND2XL U5838 ( .A(N5999), .B(n3694), .Z(n2673) );
  CANR2XL U5839 ( .A(mem_data1[841]), .B(n3898), .C(N9121), .D(n3662), .Z(
        n2672) );
  CANR2XL U5840 ( .A(N2916), .B(n3575), .C(n3611), .D(N7439), .Z(n2677) );
  CND2XL U5841 ( .A(N5998), .B(n3691), .Z(n2676) );
  CANR2XL U5842 ( .A(mem_data1[840]), .B(n3898), .C(N9120), .D(n3662), .Z(
        n2675) );
  CANR2XL U5843 ( .A(N2915), .B(n3575), .C(n3611), .D(N7440), .Z(n2680) );
  CND2XL U5844 ( .A(N5997), .B(n3696), .Z(n2679) );
  CANR2XL U5845 ( .A(mem_data1[839]), .B(n3898), .C(N9119), .D(n3662), .Z(
        n2678) );
  CANR2XL U5846 ( .A(N2914), .B(n3575), .C(n3611), .D(N7441), .Z(n2683) );
  CND2XL U5847 ( .A(N5996), .B(n3695), .Z(n2682) );
  CANR2XL U5848 ( .A(mem_data1[838]), .B(n3898), .C(N9118), .D(n3662), .Z(
        n2681) );
  CANR2XL U5849 ( .A(N2913), .B(n3575), .C(n3611), .D(N7442), .Z(n2686) );
  CND2XL U5850 ( .A(N5995), .B(n3690), .Z(n2685) );
  CANR2XL U5851 ( .A(mem_data1[837]), .B(n3898), .C(N9117), .D(n3662), .Z(
        n2684) );
  CANR2XL U5852 ( .A(N2912), .B(n3577), .C(n3611), .D(N7443), .Z(n2689) );
  CND2XL U5853 ( .A(N5994), .B(n3694), .Z(n2688) );
  CANR2XL U5854 ( .A(mem_data1[836]), .B(n3898), .C(N9116), .D(n3662), .Z(
        n2687) );
  CANR2XL U5855 ( .A(N2911), .B(n3577), .C(n3611), .D(N7444), .Z(n2692) );
  CND2XL U5856 ( .A(N5993), .B(n3691), .Z(n2691) );
  CANR2XL U5857 ( .A(mem_data1[835]), .B(n3898), .C(N9115), .D(n3662), .Z(
        n2690) );
  CANR2XL U5858 ( .A(N2910), .B(n3577), .C(n3611), .D(N7445), .Z(n2695) );
  CND2XL U5859 ( .A(N5992), .B(n3696), .Z(n2694) );
  CANR2XL U5860 ( .A(mem_data1[834]), .B(n3898), .C(N9114), .D(n3662), .Z(
        n2693) );
  CANR2XL U5861 ( .A(N2909), .B(n3577), .C(n3611), .D(N7446), .Z(n2698) );
  CND2XL U5862 ( .A(N5991), .B(n3695), .Z(n2697) );
  CANR2XL U5863 ( .A(mem_data1[833]), .B(n3898), .C(N9113), .D(n3662), .Z(
        n2696) );
  CANR2XL U5864 ( .A(N2883), .B(n3578), .C(n3612), .D(N7472), .Z(n2776) );
  CND2XL U5865 ( .A(N5965), .B(n3690), .Z(n2775) );
  CANR2XL U5866 ( .A(mem_data1[807]), .B(n3898), .C(N9087), .D(n3661), .Z(
        n2774) );
  CANR2XL U5867 ( .A(N2882), .B(n3574), .C(n3610), .D(N7473), .Z(n2779) );
  CND2XL U5868 ( .A(N5964), .B(n3694), .Z(n2778) );
  CANR2XL U5869 ( .A(mem_data1[806]), .B(n3898), .C(N9086), .D(n3661), .Z(
        n2777) );
  CANR2XL U5870 ( .A(N2763), .B(n3599), .C(n3632), .D(N7592), .Z(n3136) );
  CND2XL U5871 ( .A(N5845), .B(n3691), .Z(n3135) );
  CANR2XL U5872 ( .A(mem_data1[687]), .B(n3898), .C(N8967), .D(n3665), .Z(
        n3134) );
  CANR2XL U5873 ( .A(N2762), .B(n3599), .C(n3632), .D(N7593), .Z(n3139) );
  CND2XL U5874 ( .A(N5844), .B(n3691), .Z(n3138) );
  CANR2XL U5875 ( .A(mem_data1[686]), .B(n3898), .C(N8966), .D(n3665), .Z(
        n3137) );
  CANR2XL U5876 ( .A(N2761), .B(n3599), .C(n3632), .D(N7594), .Z(n3142) );
  CND2XL U5877 ( .A(N5843), .B(n3698), .Z(n3141) );
  CANR2XL U5878 ( .A(mem_data1[685]), .B(n3898), .C(N8965), .D(n3665), .Z(
        n3140) );
  CANR2XL U5879 ( .A(N2760), .B(n3599), .C(n3632), .D(N7595), .Z(n3145) );
  CND2XL U5880 ( .A(N5842), .B(n3694), .Z(n3144) );
  CANR2XL U5881 ( .A(mem_data1[684]), .B(n3898), .C(N8964), .D(n3665), .Z(
        n3143) );
  CANR2XL U5882 ( .A(N2759), .B(n3599), .C(n3632), .D(N7596), .Z(n3148) );
  CND2XL U5883 ( .A(N5841), .B(n3686), .Z(n3147) );
  CANR2XL U5884 ( .A(mem_data1[683]), .B(n3898), .C(N8963), .D(n3665), .Z(
        n3146) );
  CANR2XL U5885 ( .A(N2758), .B(n3598), .C(n3632), .D(N7597), .Z(n3151) );
  CND2XL U5886 ( .A(N5840), .B(n3698), .Z(n3150) );
  CANR2XL U5887 ( .A(mem_data1[682]), .B(n3898), .C(N8962), .D(n3665), .Z(
        n3149) );
  CANR2XL U5888 ( .A(N2757), .B(n3598), .C(n3632), .D(N7598), .Z(n3154) );
  CND2XL U5889 ( .A(N5839), .B(n3683), .Z(n3153) );
  CANR2XL U5890 ( .A(mem_data1[681]), .B(n3898), .C(N8961), .D(n3665), .Z(
        n3152) );
  CANR2XL U5891 ( .A(N2756), .B(n3598), .C(n3632), .D(N7599), .Z(n3157) );
  CND2XL U5892 ( .A(N5838), .B(n3691), .Z(n3156) );
  CANR2XL U5893 ( .A(mem_data1[680]), .B(n3898), .C(N8960), .D(n3665), .Z(
        n3155) );
  CANR2XL U5894 ( .A(N2755), .B(n3600), .C(n3632), .D(N7600), .Z(n3160) );
  CND2XL U5895 ( .A(N5837), .B(n3689), .Z(n3159) );
  CANR2XL U5896 ( .A(mem_data1[679]), .B(n3898), .C(N8959), .D(n3665), .Z(
        n3158) );
  CANR2XL U5897 ( .A(N2754), .B(n3597), .C(n3630), .D(N7601), .Z(n3163) );
  CND2XL U5898 ( .A(N5836), .B(n3689), .Z(n3162) );
  CANR2XL U5899 ( .A(mem_data1[678]), .B(n3898), .C(N8958), .D(n3665), .Z(
        n3161) );
  CANR2XL U5900 ( .A(N2753), .B(n3591), .C(n3635), .D(N7602), .Z(n3166) );
  CND2XL U5901 ( .A(N5835), .B(n3690), .Z(n3165) );
  CANR2XL U5902 ( .A(mem_data1[677]), .B(n3898), .C(N8957), .D(n3665), .Z(
        n3164) );
  CANR2XL U5903 ( .A(N2751), .B(n3572), .C(n3612), .D(N7604), .Z(n78) );
  CND2XL U5904 ( .A(N5833), .B(n3687), .Z(n77) );
  CANR2XL U5905 ( .A(mem_data1[675]), .B(n3898), .C(N8955), .D(n3665), .Z(n76)
         );
  CANR2XL U5906 ( .A(N2750), .B(n3572), .C(n3608), .D(N7605), .Z(n82) );
  CND2XL U5907 ( .A(N5832), .B(n3687), .Z(n81) );
  CANR2XL U5908 ( .A(mem_data1[674]), .B(n3898), .C(N8954), .D(n3665), .Z(n80)
         );
  CANR2XL U5909 ( .A(N2749), .B(n3572), .C(n3608), .D(N7606), .Z(n85) );
  CND2XL U5910 ( .A(N5831), .B(n3687), .Z(n84) );
  CANR2XL U5911 ( .A(mem_data1[673]), .B(n3898), .C(N8953), .D(n3665), .Z(n83)
         );
  CND2XL U5912 ( .A(N5830), .B(n3687), .Z(n87) );
  CANR2XL U5913 ( .A(mem_data1[672]), .B(n3898), .C(N8952), .D(n3665), .Z(n86)
         );
  CANR2XL U5914 ( .A(N2747), .B(n3572), .C(n3608), .D(N7608), .Z(n91) );
  CND2XL U5915 ( .A(N5829), .B(n3687), .Z(n90) );
  CANR2XL U5916 ( .A(mem_data1[671]), .B(n3898), .C(N8951), .D(n3665), .Z(n89)
         );
  CANR2XL U5917 ( .A(N2746), .B(n3572), .C(n3608), .D(N7609), .Z(n94) );
  CND2XL U5918 ( .A(N5828), .B(n3687), .Z(n93) );
  CANR2XL U5919 ( .A(mem_data1[670]), .B(n3898), .C(N8950), .D(n3665), .Z(n92)
         );
  CANR2XL U5920 ( .A(N2745), .B(n3572), .C(n3607), .D(N7610), .Z(n97) );
  CND2XL U5921 ( .A(N5827), .B(n3687), .Z(n96) );
  CANR2XL U5922 ( .A(mem_data1[669]), .B(n3898), .C(N8949), .D(n3665), .Z(n95)
         );
  CANR2XL U5923 ( .A(N2744), .B(n3572), .C(n3607), .D(N7611), .Z(n100) );
  CND2XL U5924 ( .A(N5826), .B(n3687), .Z(n99) );
  CANR2XL U5925 ( .A(mem_data1[668]), .B(n3898), .C(N8948), .D(n3665), .Z(n98)
         );
  CANR2XL U5926 ( .A(N2743), .B(n3572), .C(n3607), .D(N7612), .Z(n103) );
  CND2XL U5927 ( .A(N5825), .B(n3687), .Z(n102) );
  CANR2XL U5928 ( .A(mem_data1[667]), .B(n3898), .C(N8947), .D(n3665), .Z(n101) );
  CANR2XL U5929 ( .A(N2721), .B(n3572), .C(n3608), .D(N7634), .Z(n169) );
  CND2XL U5930 ( .A(N5803), .B(n3691), .Z(n168) );
  CANR2XL U5931 ( .A(mem_data1[645]), .B(n3898), .C(N8925), .D(n3651), .Z(n167) );
  CANR2XL U5932 ( .A(N2720), .B(n3572), .C(n3608), .D(N7635), .Z(n172) );
  CND2XL U5933 ( .A(N5802), .B(n3686), .Z(n171) );
  CANR2XL U5934 ( .A(mem_data1[644]), .B(n3898), .C(N8924), .D(n3651), .Z(n170) );
  CANR2XL U5935 ( .A(N2719), .B(n3572), .C(n3608), .D(N7636), .Z(n175) );
  CND2XL U5936 ( .A(N5801), .B(n3698), .Z(n174) );
  CANR2XL U5937 ( .A(mem_data1[643]), .B(n3898), .C(N8923), .D(n3651), .Z(n173) );
  CANR2XL U5938 ( .A(N2718), .B(n3572), .C(n3608), .D(N7637), .Z(n178) );
  CANR2XL U5939 ( .A(mem_data1[642]), .B(n3898), .C(N8922), .D(n3651), .Z(n176) );
  CANR2XL U5940 ( .A(mem_data1[482]), .B(n3898), .C(n3643), .D(N8762), .Z(n656) );
  CND2XL U5941 ( .A(N5640), .B(n3694), .Z(n657) );
  CANR2XL U5942 ( .A(mem_data1[479]), .B(n3898), .C(n3643), .D(N8759), .Z(n665) );
  CND2XL U5943 ( .A(N5637), .B(n3688), .Z(n666) );
  CANR2XL U5944 ( .A(N2554), .B(n3571), .C(n3607), .D(N7801), .Z(n670) );
  CND2XL U5945 ( .A(N5636), .B(n3697), .Z(n669) );
  CANR2XL U5946 ( .A(mem_data1[478]), .B(n3898), .C(n3643), .D(N8758), .Z(n668) );
  CANR2XL U5947 ( .A(N2552), .B(n3571), .C(n3607), .D(N7803), .Z(n676) );
  CND2XL U5948 ( .A(N5634), .B(n3696), .Z(n675) );
  CANR2XL U5949 ( .A(mem_data1[476]), .B(n3898), .C(n3643), .D(N8756), .Z(n674) );
  CND2XL U5950 ( .A(N5633), .B(n3688), .Z(n678) );
  CANR2XL U5951 ( .A(N2551), .B(n3571), .C(n3607), .D(N7804), .Z(n679) );
  CANR2XL U5952 ( .A(N2550), .B(n3571), .C(n3607), .D(N7805), .Z(n682) );
  CND2XL U5953 ( .A(N5632), .B(n3687), .Z(n681) );
  CANR2XL U5954 ( .A(mem_data1[474]), .B(n3898), .C(n3643), .D(N8754), .Z(n680) );
  CND2XL U5955 ( .A(N5631), .B(n3685), .Z(n684) );
  CANR2XL U5956 ( .A(N2549), .B(n3571), .C(n3607), .D(N7806), .Z(n685) );
  CANR2XL U5957 ( .A(N2548), .B(n3571), .C(n3607), .D(N7807), .Z(n688) );
  CND2XL U5958 ( .A(N5630), .B(n3688), .Z(n687) );
  CANR2XL U5959 ( .A(mem_data1[472]), .B(n3898), .C(n3643), .D(N8752), .Z(n686) );
  CANR2XL U5960 ( .A(N2547), .B(n3571), .C(n3607), .D(N7808), .Z(n691) );
  CND2XL U5961 ( .A(N5629), .B(n3685), .Z(n690) );
  CANR2XL U5962 ( .A(mem_data1[471]), .B(n3898), .C(n3643), .D(N8751), .Z(n689) );
  CANR2XL U5963 ( .A(N2546), .B(n3571), .C(n3606), .D(N7809), .Z(n694) );
  CND2XL U5964 ( .A(N5628), .B(n3688), .Z(n693) );
  CANR2XL U5965 ( .A(mem_data1[470]), .B(n3898), .C(n3643), .D(N8750), .Z(n692) );
  CND2XL U5966 ( .A(N5627), .B(n3698), .Z(n696) );
  CANR2XL U5967 ( .A(N2545), .B(n3571), .C(n3606), .D(N7810), .Z(n697) );
  CANR2XL U5968 ( .A(N2544), .B(n3571), .C(n3606), .D(N7811), .Z(n700) );
  CND2XL U5969 ( .A(N5626), .B(n3691), .Z(n699) );
  CANR2XL U5970 ( .A(mem_data1[468]), .B(n3898), .C(n3643), .D(N8748), .Z(n698) );
  CANR2XL U5971 ( .A(N2543), .B(n3571), .C(n3607), .D(N7812), .Z(n703) );
  CND2XL U5972 ( .A(N5625), .B(n3685), .Z(n702) );
  CANR2XL U5973 ( .A(mem_data1[467]), .B(n3898), .C(n3643), .D(N8747), .Z(n701) );
  CANR2XL U5974 ( .A(N2542), .B(n3571), .C(n3606), .D(N7813), .Z(n706) );
  CND2XL U5975 ( .A(N5624), .B(n3698), .Z(n705) );
  CANR2XL U5976 ( .A(mem_data1[466]), .B(n3898), .C(n3643), .D(N8746), .Z(n704) );
  CND2XL U5977 ( .A(N5622), .B(n3686), .Z(n711) );
  CANR2XL U5978 ( .A(N2540), .B(n3571), .C(n3606), .D(N7815), .Z(n712) );
  CANR2XL U5979 ( .A(N2538), .B(n3571), .C(n3606), .D(N7817), .Z(n718) );
  CND2XL U5980 ( .A(N5620), .B(n3693), .Z(n717) );
  CANR2XL U5981 ( .A(mem_data1[462]), .B(n3898), .C(n3643), .D(N8742), .Z(n716) );
  CND2XL U5982 ( .A(N5619), .B(n3698), .Z(n720) );
  CANR2XL U5983 ( .A(N2537), .B(n3571), .C(n3606), .D(N7818), .Z(n721) );
  CND2XL U5984 ( .A(N5618), .B(n3684), .Z(n723) );
  CANR2XL U5985 ( .A(N2536), .B(n3570), .C(n3606), .D(N7819), .Z(n724) );
  CANR2XL U5986 ( .A(N2535), .B(n3571), .C(n3607), .D(N7820), .Z(n727) );
  CND2XL U5987 ( .A(N5617), .B(n3686), .Z(n726) );
  CANR2XL U5988 ( .A(mem_data1[459]), .B(n3898), .C(n3643), .D(N8739), .Z(n725) );
  CANR2XL U5989 ( .A(N2534), .B(n3570), .C(n3607), .D(N7821), .Z(n730) );
  CND2XL U5990 ( .A(N5616), .B(n3686), .Z(n729) );
  CANR2XL U5991 ( .A(mem_data1[458]), .B(n3898), .C(n3643), .D(N8738), .Z(n728) );
  CND2XL U5992 ( .A(N5615), .B(n3693), .Z(n732) );
  CANR2XL U5993 ( .A(N2533), .B(n3570), .C(n3607), .D(N7822), .Z(n733) );
  CANR2XL U5994 ( .A(N2532), .B(n3570), .C(n3607), .D(N7823), .Z(n736) );
  CND2XL U5995 ( .A(N5614), .B(n3697), .Z(n735) );
  CANR2XL U5996 ( .A(mem_data1[456]), .B(n3898), .C(n3643), .D(N8736), .Z(n734) );
  CANR2XL U5997 ( .A(N2530), .B(n3570), .C(n3607), .D(N7825), .Z(n742) );
  CND2XL U5998 ( .A(N5612), .B(n3696), .Z(n741) );
  CANR2XL U5999 ( .A(mem_data1[454]), .B(n3898), .C(n3643), .D(N8734), .Z(n740) );
  CANR2XL U6000 ( .A(N2528), .B(n3571), .C(n3607), .D(N7827), .Z(n748) );
  CND2XL U6001 ( .A(N5610), .B(n3698), .Z(n747) );
  CANR2XL U6002 ( .A(mem_data1[452]), .B(n3898), .C(n3643), .D(N8732), .Z(n746) );
  CND2XL U6003 ( .A(N5609), .B(n3689), .Z(n750) );
  CANR2XL U6004 ( .A(N2527), .B(n3571), .C(n3607), .D(N7828), .Z(n751) );
  CND2XL U6005 ( .A(N5608), .B(n3687), .Z(n753) );
  CANR2XL U6006 ( .A(N2526), .B(n3571), .C(n3607), .D(N7829), .Z(n754) );
  CANR2XL U6007 ( .A(N2524), .B(n3571), .C(n3607), .D(N7831), .Z(n760) );
  CND2XL U6008 ( .A(N5606), .B(n3694), .Z(n759) );
  CANR2XL U6009 ( .A(mem_data1[448]), .B(n3898), .C(n3642), .D(N8728), .Z(n758) );
  CANR2XL U6010 ( .A(mem_data1[447]), .B(n3898), .C(n3643), .D(N8727), .Z(n761) );
  CND2XL U6011 ( .A(N5605), .B(n3696), .Z(n762) );
  CND2XL U6012 ( .A(N5604), .B(n3698), .Z(n765) );
  CANR2XL U6013 ( .A(mem_data1[446]), .B(n3898), .C(n3679), .D(N8726), .Z(n764) );
  CANR2XL U6014 ( .A(mem_data1[443]), .B(n3898), .C(N8723), .D(n3679), .Z(n773) );
  CND2XL U6015 ( .A(N5592), .B(n3694), .Z(n801) );
  CANR2XL U6016 ( .A(N2510), .B(n3571), .C(n3607), .D(N7845), .Z(n802) );
  CND2XL U6017 ( .A(N5587), .B(n3687), .Z(n816) );
  CANR2XL U6018 ( .A(N2505), .B(n3571), .C(n3608), .D(N7850), .Z(n817) );
  CANR2XL U6019 ( .A(mem_data1[424]), .B(n3898), .C(n3642), .D(N8704), .Z(n830) );
  CND2XL U6020 ( .A(N5582), .B(n3686), .Z(n831) );
  CANR2XL U6021 ( .A(mem_data1[422]), .B(n3898), .C(n3642), .D(N8702), .Z(n836) );
  CND2XL U6022 ( .A(N5580), .B(n3698), .Z(n837) );
  CANR2XL U6023 ( .A(mem_data1[420]), .B(n3898), .C(n3642), .D(N8700), .Z(n842) );
  CND2XL U6024 ( .A(N5578), .B(n3689), .Z(n843) );
  CANR2XL U6025 ( .A(mem_data1[418]), .B(n3898), .C(n3642), .D(N8698), .Z(n848) );
  CND2XL U6026 ( .A(N5576), .B(n3689), .Z(n849) );
  CND2XL U6027 ( .A(N5575), .B(n3689), .Z(n852) );
  CANR2XL U6028 ( .A(mem_data1[417]), .B(n3898), .C(n3678), .D(N8697), .Z(n851) );
  CANR2XL U6029 ( .A(N2490), .B(n3580), .C(n3616), .D(N7865), .Z(n862) );
  CND2XL U6030 ( .A(N5572), .B(n3689), .Z(n861) );
  CANR2XL U6031 ( .A(mem_data1[414]), .B(n3898), .C(n3642), .D(N8694), .Z(n860) );
  CND2XL U6032 ( .A(N5570), .B(n3689), .Z(n867) );
  CANR2XL U6033 ( .A(N2488), .B(n3580), .C(n3616), .D(N7867), .Z(n868) );
  CND2XL U6034 ( .A(N5569), .B(n3689), .Z(n870) );
  CANR2XL U6035 ( .A(N2487), .B(n3580), .C(n3616), .D(N7868), .Z(n871) );
  CND2XL U6036 ( .A(N5568), .B(n3689), .Z(n873) );
  CANR2XL U6037 ( .A(N2486), .B(n3580), .C(n3616), .D(N7869), .Z(n874) );
  CND2XL U6038 ( .A(N5567), .B(n3689), .Z(n876) );
  CANR2XL U6039 ( .A(N2485), .B(n3581), .C(n3616), .D(N7870), .Z(n877) );
  CND2XL U6040 ( .A(N5566), .B(n3689), .Z(n879) );
  CANR2XL U6041 ( .A(N2484), .B(n3581), .C(n3616), .D(N7871), .Z(n880) );
  CND2XL U6042 ( .A(N5565), .B(n3689), .Z(n882) );
  CANR2XL U6043 ( .A(N2483), .B(n3581), .C(n3616), .D(N7872), .Z(n883) );
  CANR2XL U6044 ( .A(N2482), .B(n3581), .C(n3616), .D(N7873), .Z(n886) );
  CND2XL U6045 ( .A(N5564), .B(n3689), .Z(n885) );
  CANR2XL U6046 ( .A(mem_data1[406]), .B(n3898), .C(n3642), .D(N8686), .Z(n884) );
  CND2XL U6047 ( .A(N5563), .B(n3689), .Z(n888) );
  CANR2XL U6048 ( .A(N2481), .B(n3581), .C(n3616), .D(N7874), .Z(n889) );
  CND2XL U6049 ( .A(N5562), .B(n3689), .Z(n891) );
  CANR2XL U6050 ( .A(N2480), .B(n3581), .C(n3616), .D(N7875), .Z(n892) );
  CANR2XL U6051 ( .A(mem_data1[403]), .B(n3898), .C(n3642), .D(N8683), .Z(n893) );
  CND2XL U6052 ( .A(N5561), .B(n3689), .Z(n894) );
  CND2XL U6053 ( .A(N5560), .B(n3689), .Z(n897) );
  CANR2XL U6054 ( .A(N2478), .B(n3581), .C(n3616), .D(N7877), .Z(n898) );
  CND2XL U6055 ( .A(N5556), .B(n3687), .Z(n909) );
  CANR2XL U6056 ( .A(N2474), .B(n3581), .C(n3616), .D(N7881), .Z(n910) );
  CND2XL U6057 ( .A(N5555), .B(n3686), .Z(n912) );
  CANR2XL U6058 ( .A(N2473), .B(n3581), .C(n3616), .D(N7882), .Z(n913) );
  CND2XL U6059 ( .A(N5554), .B(n3687), .Z(n915) );
  CANR2XL U6060 ( .A(N2472), .B(n3581), .C(n3616), .D(N7883), .Z(n916) );
  CND2XL U6061 ( .A(N5551), .B(n3693), .Z(n924) );
  CANR2XL U6062 ( .A(N2469), .B(n3581), .C(n3616), .D(N7886), .Z(n925) );
  CANR2XL U6063 ( .A(N2468), .B(n3581), .C(n3617), .D(N7887), .Z(n928) );
  CND2XL U6064 ( .A(N5550), .B(n3698), .Z(n927) );
  CANR2XL U6065 ( .A(mem_data1[392]), .B(n3898), .C(n3642), .D(N8672), .Z(n926) );
  CANR2XL U6066 ( .A(N2466), .B(n3581), .C(n3617), .D(N7889), .Z(n934) );
  CND2XL U6067 ( .A(N5548), .B(n3694), .Z(n933) );
  CANR2XL U6068 ( .A(mem_data1[390]), .B(n3898), .C(n3642), .D(N8670), .Z(n932) );
  CND2XL U6069 ( .A(N5547), .B(n3694), .Z(n936) );
  CANR2XL U6070 ( .A(N2465), .B(n3581), .C(n3617), .D(N7890), .Z(n937) );
  CND2XL U6071 ( .A(N5546), .B(n3690), .Z(n939) );
  CANR2XL U6072 ( .A(N2464), .B(n3581), .C(n3617), .D(N7891), .Z(n940) );
  CND2XL U6073 ( .A(N5545), .B(n3693), .Z(n942) );
  CANR2XL U6074 ( .A(N2463), .B(n3581), .C(n3616), .D(N7892), .Z(n943) );
  CND2XL U6075 ( .A(N5544), .B(n3689), .Z(n945) );
  CANR2XL U6076 ( .A(N2462), .B(n3581), .C(n3616), .D(N7893), .Z(n946) );
  CND2XL U6077 ( .A(N5543), .B(n3693), .Z(n948) );
  CANR2XL U6078 ( .A(N2461), .B(n3581), .C(n3616), .D(N7894), .Z(n949) );
  CND2XL U6079 ( .A(N5542), .B(n3683), .Z(n951) );
  CANR2XL U6080 ( .A(mem_data1[384]), .B(n3898), .C(n3642), .D(N8664), .Z(n950) );
  CANR2XL U6081 ( .A(mem_data1[383]), .B(n3898), .C(n3642), .D(N8663), .Z(n953) );
  CND2XL U6082 ( .A(N5541), .B(n3691), .Z(n954) );
  CANR2XL U6083 ( .A(mem_data1[382]), .B(n3898), .C(n3642), .D(N8662), .Z(n956) );
  CND2XL U6084 ( .A(N5540), .B(n3692), .Z(n957) );
  CANR2XL U6085 ( .A(mem_data1[372]), .B(n3898), .C(n3642), .D(N8652), .Z(n986) );
  CND2XL U6086 ( .A(N5530), .B(n3693), .Z(n987) );
  CANR2XL U6087 ( .A(mem_data1[371]), .B(n3898), .C(n3641), .D(N8651), .Z(n989) );
  CND2XL U6088 ( .A(N5529), .B(n3691), .Z(n990) );
  CND2XL U6089 ( .A(N5526), .B(n3693), .Z(n999) );
  CANR2XL U6090 ( .A(mem_data1[368]), .B(n3898), .C(n3642), .D(N8648), .Z(n998) );
  CND2XL U6091 ( .A(N5524), .B(n3693), .Z(n1005) );
  CANR2XL U6092 ( .A(mem_data1[366]), .B(n3898), .C(n3678), .D(N8646), .Z(
        n1004) );
  CND2XL U6093 ( .A(N5508), .B(n3690), .Z(n1053) );
  CANR2XL U6094 ( .A(N2426), .B(n3582), .C(n3617), .D(N7929), .Z(n1054) );
  CND2XL U6095 ( .A(N5506), .B(n3690), .Z(n1059) );
  CANR2XL U6096 ( .A(N2424), .B(n3582), .C(n3617), .D(N7931), .Z(n1060) );
  CND2XL U6097 ( .A(N5504), .B(n3690), .Z(n1065) );
  CANR2XL U6098 ( .A(N2422), .B(n3582), .C(n3617), .D(N7933), .Z(n1066) );
  CND2XL U6099 ( .A(N5503), .B(n3690), .Z(n1068) );
  CANR2XL U6100 ( .A(N2421), .B(n3582), .C(n3617), .D(N7934), .Z(n1069) );
  CND2XL U6101 ( .A(N5502), .B(n3690), .Z(n1071) );
  CANR2XL U6102 ( .A(N2420), .B(n3582), .C(n3617), .D(N7935), .Z(n1072) );
  CND2XL U6103 ( .A(N5501), .B(n3690), .Z(n1074) );
  CANR2XL U6104 ( .A(N2419), .B(n3582), .C(n3617), .D(N7936), .Z(n1075) );
  CND2XL U6105 ( .A(N5500), .B(n3690), .Z(n1077) );
  CANR2XL U6106 ( .A(N2418), .B(n3582), .C(n3617), .D(N7937), .Z(n1078) );
  CND2XL U6107 ( .A(N5499), .B(n3690), .Z(n1080) );
  CANR2XL U6108 ( .A(N2417), .B(n3582), .C(n3617), .D(N7938), .Z(n1081) );
  CND2XL U6109 ( .A(N5498), .B(n3690), .Z(n1083) );
  CANR2XL U6110 ( .A(N2416), .B(n3582), .C(n3617), .D(N7939), .Z(n1084) );
  CANR2XL U6111 ( .A(N2414), .B(n3582), .C(n3618), .D(N7941), .Z(n1090) );
  CND2XL U6112 ( .A(N5496), .B(n3690), .Z(n1089) );
  CANR2XL U6113 ( .A(mem_data1[338]), .B(n3898), .C(n3641), .D(N8618), .Z(
        n1088) );
  CND2XL U6114 ( .A(N5495), .B(n3690), .Z(n1092) );
  CANR2XL U6115 ( .A(N2413), .B(n3582), .C(n3618), .D(N7942), .Z(n1093) );
  CANR2XL U6116 ( .A(N2412), .B(n3582), .C(n3618), .D(N7943), .Z(n1096) );
  CND2XL U6117 ( .A(N5494), .B(n3690), .Z(n1095) );
  CANR2XL U6118 ( .A(mem_data1[336]), .B(n3898), .C(n3641), .D(N8616), .Z(
        n1094) );
  CANR2XL U6119 ( .A(N2410), .B(n3583), .C(n3618), .D(N7945), .Z(n1102) );
  CND2XL U6120 ( .A(N5492), .B(n3688), .Z(n1101) );
  CANR2XL U6121 ( .A(mem_data1[334]), .B(n3898), .C(n3641), .D(N8614), .Z(
        n1100) );
  CANR2XL U6122 ( .A(N2409), .B(n3583), .C(n3617), .D(N7946), .Z(n1105) );
  CND2XL U6123 ( .A(N5491), .B(n3686), .Z(n1104) );
  CANR2XL U6124 ( .A(mem_data1[333]), .B(n3898), .C(n3641), .D(N8613), .Z(
        n1103) );
  CANR2XL U6125 ( .A(N2408), .B(n3583), .C(n3617), .D(N7947), .Z(n1108) );
  CND2XL U6126 ( .A(N5490), .B(n3683), .Z(n1107) );
  CANR2XL U6127 ( .A(mem_data1[332]), .B(n3898), .C(n3641), .D(N8612), .Z(
        n1106) );
  CANR2XL U6128 ( .A(mem_data1[331]), .B(n3898), .C(n3641), .D(N8611), .Z(
        n1109) );
  CND2XL U6129 ( .A(N5489), .B(n3696), .Z(n1110) );
  CANR2XL U6130 ( .A(N2406), .B(n3583), .C(n3617), .D(N7949), .Z(n1114) );
  CND2XL U6131 ( .A(N5488), .B(n3694), .Z(n1113) );
  CANR2XL U6132 ( .A(mem_data1[330]), .B(n3898), .C(n3641), .D(N8610), .Z(
        n1112) );
  CANR2XL U6133 ( .A(N2405), .B(n3582), .C(n3617), .D(N7950), .Z(n1117) );
  CND2XL U6134 ( .A(N5487), .B(n3686), .Z(n1116) );
  CANR2XL U6135 ( .A(mem_data1[329]), .B(n3898), .C(n3641), .D(N8609), .Z(
        n1115) );
  CANR2XL U6136 ( .A(N2404), .B(n3582), .C(n3617), .D(N7951), .Z(n1120) );
  CND2XL U6137 ( .A(N5486), .B(n3683), .Z(n1119) );
  CANR2XL U6138 ( .A(mem_data1[328]), .B(n3898), .C(n3641), .D(N8608), .Z(
        n1118) );
  CND2XL U6139 ( .A(N5484), .B(n3685), .Z(n1125) );
  CANR2XL U6140 ( .A(N2402), .B(n3582), .C(n3617), .D(N7953), .Z(n1126) );
  CND2XL U6141 ( .A(N5482), .B(n3696), .Z(n1131) );
  CANR2XL U6142 ( .A(N2400), .B(n3582), .C(n3617), .D(N7955), .Z(n1132) );
  CND2XL U6143 ( .A(N5481), .B(n3691), .Z(n1134) );
  CANR2XL U6144 ( .A(N2399), .B(n3582), .C(n3617), .D(N7956), .Z(n1135) );
  CANR2XL U6145 ( .A(N2398), .B(n3582), .C(n3617), .D(N7957), .Z(n1138) );
  CND2XL U6146 ( .A(N5480), .B(n3692), .Z(n1137) );
  CANR2XL U6147 ( .A(mem_data1[322]), .B(n3898), .C(n3641), .D(N8602), .Z(
        n1136) );
  CND2XL U6148 ( .A(N5479), .B(n3683), .Z(n1140) );
  CANR2XL U6149 ( .A(N2397), .B(n3582), .C(n3617), .D(N7958), .Z(n1141) );
  CANR2XL U6150 ( .A(mem_data1[319]), .B(n3898), .C(n3641), .D(N8599), .Z(
        n1145) );
  CND2XL U6151 ( .A(N5477), .B(n3691), .Z(n1146) );
  CANR2XL U6152 ( .A(mem_data1[318]), .B(n3898), .C(n3641), .D(N8598), .Z(
        n1148) );
  CND2XL U6153 ( .A(N5476), .B(n3685), .Z(n1149) );
  CND2XL U6154 ( .A(N5474), .B(n3688), .Z(n1155) );
  CANR2XL U6155 ( .A(mem_data1[316]), .B(n3898), .C(n3678), .D(N8596), .Z(
        n1154) );
  CND2XL U6156 ( .A(N5472), .B(n3697), .Z(n1161) );
  CANR2XL U6157 ( .A(mem_data1[314]), .B(n3898), .C(n3678), .D(N8594), .Z(
        n1160) );
  CANR2XL U6158 ( .A(mem_data1[312]), .B(n3898), .C(n3641), .D(N8592), .Z(
        n1166) );
  CND2XL U6159 ( .A(N5470), .B(n3694), .Z(n1167) );
  CANR2XL U6160 ( .A(N2387), .B(n3582), .C(n3606), .D(N7968), .Z(n1171) );
  CND2XL U6161 ( .A(N5469), .B(n3690), .Z(n1170) );
  CANR2XL U6162 ( .A(mem_data1[311]), .B(n3898), .C(n3641), .D(N8591), .Z(
        n1169) );
  CANR2XL U6163 ( .A(mem_data1[310]), .B(n3898), .C(n3641), .D(N8590), .Z(
        n1172) );
  CND2XL U6164 ( .A(N5468), .B(n3690), .Z(n1173) );
  CANR2XL U6165 ( .A(mem_data1[308]), .B(n3898), .C(n3641), .D(N8588), .Z(
        n1178) );
  CND2XL U6166 ( .A(N5466), .B(n3693), .Z(n1179) );
  CANR2XL U6167 ( .A(mem_data1[307]), .B(n3898), .C(n3641), .D(N8587), .Z(
        n1181) );
  CND2XL U6168 ( .A(N5465), .B(n3686), .Z(n1182) );
  CND2XL U6169 ( .A(N5462), .B(n3691), .Z(n1191) );
  CANR2XL U6170 ( .A(N2380), .B(n3583), .C(n3618), .D(N7975), .Z(n1192) );
  CND2XL U6171 ( .A(N5459), .B(n3687), .Z(n1200) );
  CANR2XL U6172 ( .A(N2377), .B(n3583), .C(n3618), .D(N7978), .Z(n1201) );
  CANR2XL U6173 ( .A(mem_data1[289]), .B(n3898), .C(n3641), .D(N8569), .Z(
        n1235) );
  CND2XL U6174 ( .A(N5447), .B(n3687), .Z(n1236) );
  CANR2XL U6175 ( .A(N2362), .B(n3585), .C(n3620), .D(N7993), .Z(n1246) );
  CND2XL U6176 ( .A(N5441), .B(n3693), .Z(n1254) );
  CANR2XL U6177 ( .A(N2359), .B(n3585), .C(n3620), .D(N7996), .Z(n1255) );
  CND2XL U6178 ( .A(N5440), .B(n3698), .Z(n1257) );
  CANR2XL U6179 ( .A(N2358), .B(n3585), .C(n3620), .D(N7997), .Z(n1258) );
  CND2XL U6180 ( .A(N5437), .B(n3688), .Z(n1266) );
  CANR2XL U6181 ( .A(N2355), .B(n3585), .C(n3620), .D(N8000), .Z(n1267) );
  CND2XL U6182 ( .A(N5436), .B(n3693), .Z(n1269) );
  CANR2XL U6183 ( .A(N2354), .B(n3585), .C(n3620), .D(N8001), .Z(n1270) );
  CND2XL U6184 ( .A(N5435), .B(n3686), .Z(n1272) );
  CANR2XL U6185 ( .A(N2353), .B(n3586), .C(n3620), .D(N8002), .Z(n1273) );
  CND2XL U6186 ( .A(N5431), .B(n3698), .Z(n1284) );
  CANR2XL U6187 ( .A(N2349), .B(n3586), .C(n3621), .D(N8006), .Z(n1285) );
  CANR2XL U6188 ( .A(N2340), .B(n3586), .C(n3621), .D(N8015), .Z(n1312) );
  CND2XL U6189 ( .A(N5422), .B(n3686), .Z(n1311) );
  CANR2XL U6190 ( .A(mem_data1[264]), .B(n3898), .C(n3642), .D(N8544), .Z(
        n1310) );
  CANR2XL U6191 ( .A(mem_data1[263]), .B(n3898), .C(n3644), .D(N8543), .Z(
        n1313) );
  CND2XL U6192 ( .A(N5421), .B(n3687), .Z(n1314) );
  CANR2XL U6193 ( .A(N2336), .B(n3586), .C(n3621), .D(N8019), .Z(n1324) );
  CND2XL U6194 ( .A(N5418), .B(n3688), .Z(n1323) );
  CANR2XL U6195 ( .A(mem_data1[260]), .B(n3898), .C(n3642), .D(N8540), .Z(
        n1322) );
  CND2XL U6196 ( .A(N5417), .B(n3696), .Z(n1326) );
  CANR2XL U6197 ( .A(N2335), .B(n3586), .C(n3621), .D(N8020), .Z(n1327) );
  CANR2XL U6198 ( .A(N2334), .B(n3586), .C(n3621), .D(N8021), .Z(n1330) );
  CND2XL U6199 ( .A(N5416), .B(n3696), .Z(n1329) );
  CANR2XL U6200 ( .A(mem_data1[258]), .B(n3898), .C(n3642), .D(N8538), .Z(
        n1328) );
  CND2XL U6201 ( .A(N5415), .B(n3694), .Z(n1332) );
  CANR2XL U6202 ( .A(N2333), .B(n3586), .C(n3621), .D(N8022), .Z(n1333) );
  CANR2XL U6203 ( .A(mem_data1[255]), .B(n3898), .C(n3642), .D(N8535), .Z(
        n1337) );
  CND2XL U6204 ( .A(N5413), .B(n3688), .Z(n1338) );
  CANR2XL U6205 ( .A(mem_data1[254]), .B(n3898), .C(n3643), .D(N8534), .Z(
        n1340) );
  CND2XL U6206 ( .A(N5412), .B(n3683), .Z(n1341) );
  CND2XL U6207 ( .A(N5400), .B(n3694), .Z(n1377) );
  CANR2XL U6208 ( .A(N2318), .B(n3587), .C(n3622), .D(N8037), .Z(n1378) );
  CANR2XL U6209 ( .A(mem_data1[241]), .B(n3898), .C(N8521), .D(n3648), .Z(
        n1379) );
  CND2XL U6210 ( .A(N5399), .B(n3693), .Z(n1380) );
  CANR2XL U6211 ( .A(N2316), .B(n3587), .C(n3622), .D(N8039), .Z(n1384) );
  CND2XL U6212 ( .A(N5398), .B(n3696), .Z(n1383) );
  CANR2XL U6213 ( .A(mem_data1[240]), .B(n3898), .C(N8520), .D(n3648), .Z(
        n1382) );
  CANR2XL U6214 ( .A(mem_data1[239]), .B(n3898), .C(N8519), .D(n3648), .Z(
        n1385) );
  CND2XL U6215 ( .A(N5397), .B(n3689), .Z(n1386) );
  CANR2XL U6216 ( .A(N2313), .B(n3587), .C(n3622), .D(N8042), .Z(n1393) );
  CND2XL U6217 ( .A(N5395), .B(n3698), .Z(n1392) );
  CANR2XL U6218 ( .A(mem_data1[237]), .B(n3898), .C(N8517), .D(n3648), .Z(
        n1391) );
  CANR2XL U6219 ( .A(N2312), .B(n3587), .C(n3622), .D(N8043), .Z(n1396) );
  CND2XL U6220 ( .A(N5394), .B(n3684), .Z(n1395) );
  CANR2XL U6221 ( .A(mem_data1[236]), .B(n3898), .C(N8516), .D(n3648), .Z(
        n1394) );
  CANR2XL U6222 ( .A(N2311), .B(n3587), .C(n3622), .D(N8044), .Z(n1399) );
  CND2XL U6223 ( .A(N5393), .B(n3692), .Z(n1398) );
  CANR2XL U6224 ( .A(mem_data1[235]), .B(n3898), .C(N8515), .D(n3648), .Z(
        n1397) );
  CND2XL U6225 ( .A(N5392), .B(n3686), .Z(n1401) );
  CANR2XL U6226 ( .A(N2310), .B(n3587), .C(n3622), .D(N8045), .Z(n1402) );
  CANR2XL U6227 ( .A(N2309), .B(n3587), .C(n3622), .D(N8046), .Z(n1405) );
  CND2XL U6228 ( .A(N5391), .B(n3687), .Z(n1404) );
  CANR2XL U6229 ( .A(mem_data1[233]), .B(n3898), .C(N8513), .D(n3648), .Z(
        n1403) );
  CANR2XL U6230 ( .A(mem_data1[232]), .B(n3898), .C(N8512), .D(n3648), .Z(
        n1406) );
  CND2XL U6231 ( .A(N5390), .B(n3689), .Z(n1407) );
  CANR2XL U6232 ( .A(mem_data1[231]), .B(n3898), .C(N8511), .D(n3648), .Z(
        n1409) );
  CND2XL U6233 ( .A(N5389), .B(n3696), .Z(n1410) );
  CANR2XL U6234 ( .A(mem_data1[229]), .B(n3898), .C(N8509), .D(n3648), .Z(
        n1415) );
  CND2XL U6235 ( .A(N5387), .B(n3697), .Z(n1416) );
  CND2XL U6236 ( .A(N5386), .B(n3697), .Z(n1419) );
  CANR2XL U6237 ( .A(N2304), .B(n3586), .C(n3622), .D(N8051), .Z(n1420) );
  CANR2XL U6238 ( .A(mem_data1[227]), .B(n3898), .C(N8507), .D(n3648), .Z(
        n1421) );
  CND2XL U6239 ( .A(N5385), .B(n3689), .Z(n1422) );
  CANR2XL U6240 ( .A(N2302), .B(n3579), .C(n3621), .D(N8053), .Z(n1426) );
  CND2XL U6241 ( .A(N5384), .B(n3686), .Z(n1425) );
  CANR2XL U6242 ( .A(mem_data1[226]), .B(n3898), .C(N8506), .D(n3648), .Z(
        n1424) );
  CANR2XL U6243 ( .A(N2301), .B(n3579), .C(n3621), .D(N8054), .Z(n1429) );
  CND2XL U6244 ( .A(N5383), .B(n3698), .Z(n1428) );
  CANR2XL U6245 ( .A(mem_data1[225]), .B(n3898), .C(N8505), .D(n3648), .Z(
        n1427) );
  CANR2XL U6246 ( .A(N2300), .B(n3579), .C(n3621), .D(N8055), .Z(n1432) );
  CND2XL U6247 ( .A(N5382), .B(n3693), .Z(n1431) );
  CANR2XL U6248 ( .A(mem_data1[224]), .B(n3898), .C(N8504), .D(n3648), .Z(
        n1430) );
  CANR2XL U6249 ( .A(N2299), .B(n3579), .C(n3621), .D(N8056), .Z(n1435) );
  CND2XL U6250 ( .A(N5381), .B(n3691), .Z(n1434) );
  CANR2XL U6251 ( .A(mem_data1[223]), .B(n3898), .C(N8503), .D(n3648), .Z(
        n1433) );
  CND2XL U6252 ( .A(N5378), .B(n3696), .Z(n1443) );
  CANR2XL U6253 ( .A(N2296), .B(n3579), .C(n3621), .D(N8059), .Z(n1444) );
  CANR2XL U6254 ( .A(N2295), .B(n3579), .C(n3621), .D(N8060), .Z(n1447) );
  CND2XL U6255 ( .A(N5377), .B(n3686), .Z(n1446) );
  CANR2XL U6256 ( .A(mem_data1[219]), .B(n3898), .C(N8499), .D(n3649), .Z(
        n1445) );
  CANR2XL U6257 ( .A(N2294), .B(n3579), .C(n3621), .D(N8061), .Z(n1450) );
  CND2XL U6258 ( .A(N5376), .B(n3692), .Z(n1449) );
  CANR2XL U6259 ( .A(mem_data1[218]), .B(n3898), .C(N8498), .D(n3649), .Z(
        n1448) );
  CANR2XL U6260 ( .A(N2293), .B(n3579), .C(n3615), .D(N8062), .Z(n1453) );
  CND2XL U6261 ( .A(N5375), .B(n3694), .Z(n1452) );
  CANR2XL U6262 ( .A(mem_data1[217]), .B(n3898), .C(N8497), .D(n3649), .Z(
        n1451) );
  CANR2XL U6263 ( .A(N2292), .B(n3578), .C(n3615), .D(N8063), .Z(n1456) );
  CND2XL U6264 ( .A(N5374), .B(n3685), .Z(n1455) );
  CANR2XL U6265 ( .A(mem_data1[216]), .B(n3898), .C(N8496), .D(n3649), .Z(
        n1454) );
  CANR2XL U6266 ( .A(N2291), .B(n3578), .C(n3615), .D(N8064), .Z(n1459) );
  CND2XL U6267 ( .A(N5373), .B(n3696), .Z(n1458) );
  CANR2XL U6268 ( .A(mem_data1[215]), .B(n3898), .C(N8495), .D(n3649), .Z(
        n1457) );
  CANR2XL U6269 ( .A(N2290), .B(n3578), .C(n3615), .D(N8065), .Z(n1462) );
  CND2XL U6270 ( .A(N5372), .B(n3690), .Z(n1461) );
  CANR2XL U6271 ( .A(mem_data1[214]), .B(n3898), .C(N8494), .D(n3649), .Z(
        n1460) );
  CANR2XL U6272 ( .A(N2289), .B(n3581), .C(n3615), .D(N8066), .Z(n1465) );
  CND2XL U6273 ( .A(N5371), .B(n3697), .Z(n1464) );
  CANR2XL U6274 ( .A(mem_data1[213]), .B(n3898), .C(N8493), .D(n3649), .Z(
        n1463) );
  CANR2XL U6275 ( .A(N2288), .B(n3587), .C(n3614), .D(N8067), .Z(n1468) );
  CND2XL U6276 ( .A(N5370), .B(n3694), .Z(n1467) );
  CANR2XL U6277 ( .A(mem_data1[212]), .B(n3898), .C(N8492), .D(n3649), .Z(
        n1466) );
  CANR2XL U6278 ( .A(N2287), .B(n3587), .C(n3614), .D(N8068), .Z(n1471) );
  CND2XL U6279 ( .A(N5369), .B(n3685), .Z(n1470) );
  CANR2XL U6280 ( .A(mem_data1[211]), .B(n3898), .C(N8491), .D(n3649), .Z(
        n1469) );
  CANR2XL U6281 ( .A(N2286), .B(n3587), .C(n3614), .D(N8069), .Z(n1474) );
  CND2XL U6282 ( .A(N5368), .B(n3696), .Z(n1473) );
  CANR2XL U6283 ( .A(mem_data1[210]), .B(n3898), .C(N8490), .D(n3649), .Z(
        n1472) );
  CANR2XL U6284 ( .A(N2285), .B(n3587), .C(n3614), .D(N8070), .Z(n1477) );
  CND2XL U6285 ( .A(N5367), .B(n3690), .Z(n1476) );
  CANR2XL U6286 ( .A(mem_data1[209]), .B(n3898), .C(N8489), .D(n3649), .Z(
        n1475) );
  CANR2XL U6287 ( .A(N2284), .B(n3587), .C(n3614), .D(N8071), .Z(n1480) );
  CND2XL U6288 ( .A(N5366), .B(n3689), .Z(n1479) );
  CANR2XL U6289 ( .A(mem_data1[208]), .B(n3898), .C(N8488), .D(n3649), .Z(
        n1478) );
  CANR2XL U6290 ( .A(N2283), .B(n3587), .C(n3614), .D(N8072), .Z(n1483) );
  CND2XL U6291 ( .A(N5365), .B(n3694), .Z(n1482) );
  CANR2XL U6292 ( .A(mem_data1[207]), .B(n3898), .C(N8487), .D(n3649), .Z(
        n1481) );
  CANR2XL U6293 ( .A(N2282), .B(n3587), .C(n3614), .D(N8073), .Z(n1486) );
  CND2XL U6294 ( .A(N5364), .B(n3683), .Z(n1485) );
  CANR2XL U6295 ( .A(mem_data1[206]), .B(n3898), .C(N8486), .D(n3649), .Z(
        n1484) );
  CANR2XL U6296 ( .A(N2281), .B(n3587), .C(n3614), .D(N8074), .Z(n1489) );
  CND2XL U6297 ( .A(N5363), .B(n3696), .Z(n1488) );
  CANR2XL U6298 ( .A(mem_data1[205]), .B(n3898), .C(N8485), .D(n3648), .Z(
        n1487) );
  CANR2XL U6299 ( .A(N2280), .B(n3587), .C(n3614), .D(N8075), .Z(n1492) );
  CND2XL U6300 ( .A(N5362), .B(n3690), .Z(n1491) );
  CANR2XL U6301 ( .A(mem_data1[204]), .B(n3898), .C(N8484), .D(n3648), .Z(
        n1490) );
  CANR2XL U6302 ( .A(N2279), .B(n3580), .C(n3614), .D(N8076), .Z(n1495) );
  CND2XL U6303 ( .A(N5361), .B(n3685), .Z(n1494) );
  CANR2XL U6304 ( .A(mem_data1[203]), .B(n3898), .C(N8483), .D(n3648), .Z(
        n1493) );
  CANR2XL U6305 ( .A(N2278), .B(n3580), .C(n3614), .D(N8077), .Z(n1498) );
  CND2XL U6306 ( .A(N5360), .B(n3694), .Z(n1497) );
  CANR2XL U6307 ( .A(mem_data1[202]), .B(n3898), .C(N8482), .D(n3648), .Z(
        n1496) );
  CANR2XL U6308 ( .A(N2277), .B(n3580), .C(n3614), .D(N8078), .Z(n1501) );
  CND2XL U6309 ( .A(N5359), .B(n3689), .Z(n1500) );
  CANR2XL U6310 ( .A(mem_data1[201]), .B(n3898), .C(N8481), .D(n3648), .Z(
        n1499) );
  CANR2XL U6311 ( .A(N2276), .B(n3580), .C(n3614), .D(N8079), .Z(n1504) );
  CND2XL U6312 ( .A(N5358), .B(n3696), .Z(n1503) );
  CANR2XL U6313 ( .A(mem_data1[200]), .B(n3898), .C(N8480), .D(n3648), .Z(
        n1502) );
  CANR2XL U6314 ( .A(N2274), .B(n3580), .C(n3614), .D(N8081), .Z(n1510) );
  CND2XL U6315 ( .A(N5356), .B(n3694), .Z(n1509) );
  CANR2XL U6316 ( .A(mem_data1[198]), .B(n3898), .C(N8478), .D(n3650), .Z(
        n1508) );
  CANR2XL U6317 ( .A(N2273), .B(n3580), .C(n3614), .D(N8082), .Z(n1513) );
  CND2XL U6318 ( .A(N5355), .B(n3694), .Z(n1512) );
  CANR2XL U6319 ( .A(mem_data1[197]), .B(n3898), .C(N8477), .D(n3650), .Z(
        n1511) );
  CANR2XL U6320 ( .A(N2272), .B(n3580), .C(n3614), .D(N8083), .Z(n1516) );
  CND2XL U6321 ( .A(N5354), .B(n3694), .Z(n1515) );
  CANR2XL U6322 ( .A(mem_data1[196]), .B(n3898), .C(N8476), .D(n3650), .Z(
        n1514) );
  CANR2XL U6323 ( .A(N2271), .B(n3579), .C(n3614), .D(N8084), .Z(n1519) );
  CND2XL U6324 ( .A(N5353), .B(n3694), .Z(n1518) );
  CANR2XL U6325 ( .A(mem_data1[195]), .B(n3898), .C(N8475), .D(n3650), .Z(
        n1517) );
  CANR2XL U6326 ( .A(N2270), .B(n3579), .C(n3614), .D(N8085), .Z(n1522) );
  CND2XL U6327 ( .A(N5352), .B(n3694), .Z(n1521) );
  CANR2XL U6328 ( .A(mem_data1[194]), .B(n3898), .C(N8474), .D(n3650), .Z(
        n1520) );
  CANR2XL U6329 ( .A(N2269), .B(n3579), .C(n3614), .D(N8086), .Z(n1525) );
  CND2XL U6330 ( .A(N5351), .B(n3694), .Z(n1524) );
  CANR2XL U6331 ( .A(mem_data1[193]), .B(n3898), .C(N8473), .D(n3649), .Z(
        n1523) );
  CANR2XL U6332 ( .A(N2268), .B(n3579), .C(n3614), .D(N8087), .Z(n1528) );
  CND2XL U6333 ( .A(N5350), .B(n3694), .Z(n1527) );
  CANR2XL U6334 ( .A(mem_data1[192]), .B(n3898), .C(N8472), .D(n3649), .Z(
        n1526) );
  CANR2XL U6335 ( .A(N2267), .B(n3579), .C(n3616), .D(N8088), .Z(n1531) );
  CND2XL U6336 ( .A(N5349), .B(n3694), .Z(n1530) );
  CANR2XL U6337 ( .A(mem_data1[191]), .B(n3898), .C(N8471), .D(n3649), .Z(
        n1529) );
  CANR2XL U6338 ( .A(mem_data1[190]), .B(n3898), .C(N8470), .D(n3649), .Z(
        n1532) );
  CND2XL U6339 ( .A(N5348), .B(n3694), .Z(n1533) );
  CANR2XL U6340 ( .A(N2264), .B(n3579), .C(n3616), .D(N8091), .Z(n1540) );
  CND2XL U6341 ( .A(N5346), .B(n3694), .Z(n1539) );
  CANR2XL U6342 ( .A(mem_data1[188]), .B(n3898), .C(n3644), .D(N8468), .Z(
        n1538) );
  CND2XL U6343 ( .A(N5345), .B(n3694), .Z(n1542) );
  CANR2XL U6344 ( .A(N2263), .B(n3579), .C(n3615), .D(N8092), .Z(n1543) );
  CND2XL U6345 ( .A(N5344), .B(n3694), .Z(n1545) );
  CANR2XL U6346 ( .A(N2262), .B(n3579), .C(n3615), .D(N8093), .Z(n1546) );
  CND2XL U6347 ( .A(N5343), .B(n3694), .Z(n1548) );
  CANR2XL U6348 ( .A(N2261), .B(n3579), .C(n3615), .D(N8094), .Z(n1549) );
  CANR2XL U6349 ( .A(N2260), .B(n3579), .C(n3615), .D(N8095), .Z(n1552) );
  CND2XL U6350 ( .A(N5342), .B(n3694), .Z(n1551) );
  CANR2XL U6351 ( .A(mem_data1[184]), .B(n3898), .C(N8464), .D(n3650), .Z(
        n1550) );
  CND2XL U6352 ( .A(N5341), .B(n3688), .Z(n1554) );
  CANR2XL U6353 ( .A(N2259), .B(n3579), .C(n3615), .D(N8096), .Z(n1555) );
  CND2XL U6354 ( .A(N5340), .B(n3692), .Z(n1557) );
  CANR2XL U6355 ( .A(N2258), .B(n3579), .C(n3615), .D(N8097), .Z(n1558) );
  CND2XL U6356 ( .A(N5339), .B(n3691), .Z(n1560) );
  CANR2XL U6357 ( .A(N2257), .B(n3579), .C(n3615), .D(N8098), .Z(n1561) );
  CANR2XL U6358 ( .A(N2256), .B(n3579), .C(n3615), .D(N8099), .Z(n1564) );
  CND2XL U6359 ( .A(N5338), .B(n3693), .Z(n1563) );
  CANR2XL U6360 ( .A(mem_data1[180]), .B(n3898), .C(N8460), .D(n3649), .Z(
        n1562) );
  CANR2XL U6361 ( .A(N2255), .B(n3579), .C(n3615), .D(N8100), .Z(n1567) );
  CND2XL U6362 ( .A(N5337), .B(n3685), .Z(n1566) );
  CANR2XL U6363 ( .A(mem_data1[179]), .B(n3898), .C(N8459), .D(n3649), .Z(
        n1565) );
  CANR2XL U6364 ( .A(N2254), .B(n3581), .C(n3615), .D(N8101), .Z(n1570) );
  CND2XL U6365 ( .A(N5336), .B(n3691), .Z(n1569) );
  CANR2XL U6366 ( .A(mem_data1[178]), .B(n3898), .C(N8458), .D(n3649), .Z(
        n1568) );
  CANR2XL U6367 ( .A(N2253), .B(n3581), .C(n3615), .D(N8102), .Z(n1573) );
  CND2XL U6368 ( .A(N5335), .B(n3695), .Z(n1572) );
  CANR2XL U6369 ( .A(mem_data1[177]), .B(n3898), .C(N8457), .D(n3651), .Z(
        n1571) );
  CANR2XL U6370 ( .A(N2252), .B(n3580), .C(n3615), .D(N8103), .Z(n1576) );
  CND2XL U6371 ( .A(N5334), .B(n3695), .Z(n1575) );
  CANR2XL U6372 ( .A(mem_data1[176]), .B(n3898), .C(N8456), .D(n3651), .Z(
        n1574) );
  CANR2XL U6373 ( .A(N2251), .B(n3580), .C(n3615), .D(N8104), .Z(n1579) );
  CND2XL U6374 ( .A(N5333), .B(n3695), .Z(n1578) );
  CANR2XL U6375 ( .A(mem_data1[175]), .B(n3898), .C(N8455), .D(n3651), .Z(
        n1577) );
  CANR2XL U6376 ( .A(mem_data1[174]), .B(n3898), .C(N8454), .D(n3651), .Z(
        n1580) );
  CND2XL U6377 ( .A(N5332), .B(n3695), .Z(n1581) );
  CANR2XL U6378 ( .A(N2249), .B(n3580), .C(n3615), .D(N8106), .Z(n1585) );
  CND2XL U6379 ( .A(N5331), .B(n3695), .Z(n1584) );
  CANR2XL U6380 ( .A(mem_data1[173]), .B(n3898), .C(N8453), .D(n3651), .Z(
        n1583) );
  CANR2XL U6381 ( .A(N2248), .B(n3580), .C(n3615), .D(N8107), .Z(n1588) );
  CND2XL U6382 ( .A(N5330), .B(n3695), .Z(n1587) );
  CANR2XL U6383 ( .A(mem_data1[172]), .B(n3898), .C(N8452), .D(n3651), .Z(
        n1586) );
  CANR2XL U6384 ( .A(N2247), .B(n3580), .C(n3615), .D(N8108), .Z(n1591) );
  CND2XL U6385 ( .A(N5329), .B(n3695), .Z(n1590) );
  CANR2XL U6386 ( .A(mem_data1[171]), .B(n3898), .C(N8451), .D(n3650), .Z(
        n1589) );
  CANR2XL U6387 ( .A(N2246), .B(n3580), .C(n3615), .D(N8109), .Z(n1594) );
  CND2XL U6388 ( .A(N5328), .B(n3695), .Z(n1593) );
  CANR2XL U6389 ( .A(mem_data1[170]), .B(n3898), .C(N8450), .D(n3650), .Z(
        n1592) );
  CANR2XL U6390 ( .A(N2245), .B(n3580), .C(n3615), .D(N8110), .Z(n1597) );
  CND2XL U6391 ( .A(N5327), .B(n3695), .Z(n1596) );
  CANR2XL U6392 ( .A(mem_data1[169]), .B(n3898), .C(N8449), .D(n3650), .Z(
        n1595) );
  CANR2XL U6393 ( .A(N2244), .B(n3580), .C(n3615), .D(N8111), .Z(n1600) );
  CND2XL U6394 ( .A(N5326), .B(n3695), .Z(n1599) );
  CANR2XL U6395 ( .A(mem_data1[168]), .B(n3898), .C(N8448), .D(n3650), .Z(
        n1598) );
  CANR2XL U6396 ( .A(N2243), .B(n3580), .C(n3615), .D(N8112), .Z(n1603) );
  CND2XL U6397 ( .A(N5325), .B(n3695), .Z(n1602) );
  CANR2XL U6398 ( .A(mem_data1[167]), .B(n3898), .C(N8447), .D(n3651), .Z(
        n1601) );
  CANR2XL U6399 ( .A(N2242), .B(n3580), .C(n3615), .D(N8113), .Z(n1606) );
  CND2XL U6400 ( .A(N5324), .B(n3695), .Z(n1605) );
  CANR2XL U6401 ( .A(mem_data1[166]), .B(n3898), .C(N8446), .D(n3650), .Z(
        n1604) );
  CANR2XL U6402 ( .A(N2241), .B(n3580), .C(n3615), .D(N8114), .Z(n1609) );
  CND2XL U6403 ( .A(N5323), .B(n3695), .Z(n1608) );
  CANR2XL U6404 ( .A(mem_data1[165]), .B(n3898), .C(N8445), .D(n3650), .Z(
        n1607) );
  CANR2XL U6405 ( .A(N2240), .B(n3581), .C(n3616), .D(N8115), .Z(n1612) );
  CND2XL U6406 ( .A(N5322), .B(n3695), .Z(n1611) );
  CANR2XL U6407 ( .A(mem_data1[164]), .B(n3898), .C(N8444), .D(n3650), .Z(
        n1610) );
  CANR2XL U6408 ( .A(mem_data1[163]), .B(n3898), .C(N8443), .D(n3650), .Z(
        n1613) );
  CND2XL U6409 ( .A(N5321), .B(n3695), .Z(n1614) );
  CANR2XL U6410 ( .A(N2237), .B(n3580), .C(n3616), .D(N8118), .Z(n1621) );
  CND2XL U6411 ( .A(N5319), .B(n3694), .Z(n1620) );
  CANR2XL U6412 ( .A(mem_data1[161]), .B(n3898), .C(N8441), .D(n3650), .Z(
        n1619) );
  CANR2XL U6413 ( .A(N2236), .B(n3579), .C(n3621), .D(N8119), .Z(n1624) );
  CND2XL U6414 ( .A(N5318), .B(n3694), .Z(n1623) );
  CANR2XL U6415 ( .A(mem_data1[160]), .B(n3898), .C(N8440), .D(n3650), .Z(
        n1622) );
  CANR2XL U6416 ( .A(N2235), .B(n3585), .C(n3620), .D(N8120), .Z(n1627) );
  CND2XL U6417 ( .A(N5317), .B(n3694), .Z(n1626) );
  CANR2XL U6418 ( .A(mem_data1[159]), .B(n3898), .C(N8439), .D(n3650), .Z(
        n1625) );
  CANR2XL U6419 ( .A(mem_data1[158]), .B(n3898), .C(N8438), .D(n3650), .Z(
        n1628) );
  CND2XL U6420 ( .A(N5316), .B(n3694), .Z(n1629) );
  CANR2XL U6421 ( .A(N2233), .B(n3596), .C(n3622), .D(N8122), .Z(n1633) );
  CND2XL U6422 ( .A(N5315), .B(n3694), .Z(n1632) );
  CANR2XL U6423 ( .A(mem_data1[157]), .B(n3898), .C(N8437), .D(n3650), .Z(
        n1631) );
  CND2XL U6424 ( .A(N5314), .B(n3694), .Z(n1635) );
  CANR2XL U6425 ( .A(N2232), .B(n3596), .C(n3622), .D(N8123), .Z(n1636) );
  CANR2XL U6426 ( .A(N2231), .B(n3596), .C(n3622), .D(N8124), .Z(n1639) );
  CND2XL U6427 ( .A(N5313), .B(n3696), .Z(n1638) );
  CANR2XL U6428 ( .A(mem_data1[155]), .B(n3898), .C(N8435), .D(n3647), .Z(
        n1637) );
  CANR2XL U6429 ( .A(N2230), .B(n3596), .C(n3622), .D(N8125), .Z(n1642) );
  CND2XL U6430 ( .A(N5312), .B(n3696), .Z(n1641) );
  CANR2XL U6431 ( .A(mem_data1[154]), .B(n3898), .C(N8434), .D(n3647), .Z(
        n1640) );
  CANR2XL U6432 ( .A(N2229), .B(n3596), .C(n3622), .D(N8126), .Z(n1645) );
  CND2XL U6433 ( .A(N5311), .B(n3696), .Z(n1644) );
  CANR2XL U6434 ( .A(mem_data1[153]), .B(n3898), .C(N8433), .D(n3647), .Z(
        n1643) );
  CANR2XL U6435 ( .A(N2228), .B(n3596), .C(n3622), .D(N8127), .Z(n1648) );
  CND2XL U6436 ( .A(N5310), .B(n3696), .Z(n1647) );
  CANR2XL U6437 ( .A(mem_data1[152]), .B(n3898), .C(N8432), .D(n3647), .Z(
        n1646) );
  CANR2XL U6438 ( .A(N2227), .B(n3596), .C(n3622), .D(N8128), .Z(n1651) );
  CND2XL U6439 ( .A(N5309), .B(n3696), .Z(n1650) );
  CANR2XL U6440 ( .A(mem_data1[151]), .B(n3898), .C(N8431), .D(n3647), .Z(
        n1649) );
  CANR2XL U6441 ( .A(N2226), .B(n3589), .C(n3624), .D(N8129), .Z(n1654) );
  CND2XL U6442 ( .A(N5308), .B(n3696), .Z(n1653) );
  CANR2XL U6443 ( .A(mem_data1[150]), .B(n3898), .C(N8430), .D(n3647), .Z(
        n1652) );
  CANR2XL U6444 ( .A(N2225), .B(n3589), .C(n3630), .D(N8130), .Z(n1657) );
  CND2XL U6445 ( .A(N5307), .B(n3696), .Z(n1656) );
  CANR2XL U6446 ( .A(mem_data1[149]), .B(n3898), .C(N8429), .D(n3647), .Z(
        n1655) );
  CANR2XL U6447 ( .A(N2224), .B(n3589), .C(n3630), .D(N8131), .Z(n1660) );
  CND2XL U6448 ( .A(N5306), .B(n3696), .Z(n1659) );
  CANR2XL U6449 ( .A(mem_data1[148]), .B(n3898), .C(N8428), .D(n3647), .Z(
        n1658) );
  CANR2XL U6450 ( .A(N2223), .B(n3589), .C(n3630), .D(N8132), .Z(n1663) );
  CND2XL U6451 ( .A(N5305), .B(n3696), .Z(n1662) );
  CANR2XL U6452 ( .A(mem_data1[147]), .B(n3898), .C(N8427), .D(n3647), .Z(
        n1661) );
  CANR2XL U6453 ( .A(N2222), .B(n3589), .C(n3630), .D(N8133), .Z(n1666) );
  CND2XL U6454 ( .A(N5304), .B(n3696), .Z(n1665) );
  CANR2XL U6455 ( .A(mem_data1[146]), .B(n3898), .C(N8426), .D(n3650), .Z(
        n1664) );
  CANR2XL U6456 ( .A(N2221), .B(n3588), .C(n3630), .D(N8134), .Z(n1669) );
  CND2XL U6457 ( .A(N5303), .B(n3696), .Z(n1668) );
  CANR2XL U6458 ( .A(mem_data1[145]), .B(n3898), .C(N8425), .D(n3650), .Z(
        n1667) );
  CANR2XL U6459 ( .A(N2220), .B(n3588), .C(n3630), .D(N8135), .Z(n1672) );
  CND2XL U6460 ( .A(N5302), .B(n3696), .Z(n1671) );
  CANR2XL U6461 ( .A(mem_data1[144]), .B(n3898), .C(N8424), .D(n3644), .Z(
        n1670) );
  CANR2XL U6462 ( .A(N2219), .B(n3588), .C(n3630), .D(N8136), .Z(n1675) );
  CND2XL U6463 ( .A(N5301), .B(n3696), .Z(n1674) );
  CANR2XL U6464 ( .A(mem_data1[143]), .B(n3898), .C(N8423), .D(n3651), .Z(
        n1673) );
  CANR2XL U6465 ( .A(N2218), .B(n3588), .C(n3623), .D(N8137), .Z(n1678) );
  CND2XL U6466 ( .A(N5300), .B(n3696), .Z(n1677) );
  CANR2XL U6467 ( .A(mem_data1[142]), .B(n3898), .C(N8422), .D(n3651), .Z(
        n1676) );
  CANR2XL U6468 ( .A(N2217), .B(n3588), .C(n3623), .D(N8138), .Z(n1681) );
  CND2XL U6469 ( .A(N5299), .B(n3696), .Z(n1680) );
  CANR2XL U6470 ( .A(mem_data1[141]), .B(n3898), .C(N8421), .D(n3651), .Z(
        n1679) );
  CANR2XL U6471 ( .A(N2216), .B(n3588), .C(n3623), .D(N8139), .Z(n1684) );
  CND2XL U6472 ( .A(N5298), .B(n3696), .Z(n1683) );
  CANR2XL U6473 ( .A(mem_data1[140]), .B(n3898), .C(N8420), .D(n3651), .Z(
        n1682) );
  CANR2XL U6474 ( .A(N2215), .B(n3588), .C(n3623), .D(N8140), .Z(n1687) );
  CND2XL U6475 ( .A(N5297), .B(n3695), .Z(n1686) );
  CANR2XL U6476 ( .A(mem_data1[139]), .B(n3898), .C(N8419), .D(n3651), .Z(
        n1685) );
  CANR2XL U6477 ( .A(N2214), .B(n3588), .C(n3623), .D(N8141), .Z(n1690) );
  CND2XL U6478 ( .A(N5296), .B(n3695), .Z(n1689) );
  CANR2XL U6479 ( .A(mem_data1[138]), .B(n3898), .C(N8418), .D(n3651), .Z(
        n1688) );
  CANR2XL U6480 ( .A(N2213), .B(n3588), .C(n3623), .D(N8142), .Z(n1693) );
  CND2XL U6481 ( .A(N5295), .B(n3695), .Z(n1692) );
  CANR2XL U6482 ( .A(mem_data1[137]), .B(n3898), .C(N8417), .D(n3651), .Z(
        n1691) );
  CANR2XL U6483 ( .A(N2212), .B(n3588), .C(n3623), .D(N8143), .Z(n1696) );
  CND2XL U6484 ( .A(N5294), .B(n3695), .Z(n1695) );
  CANR2XL U6485 ( .A(mem_data1[136]), .B(n3898), .C(N8416), .D(n3651), .Z(
        n1694) );
  CANR2XL U6486 ( .A(N2211), .B(n3588), .C(n3623), .D(N8144), .Z(n1699) );
  CND2XL U6487 ( .A(N5293), .B(n3695), .Z(n1698) );
  CANR2XL U6488 ( .A(mem_data1[135]), .B(n3898), .C(N8415), .D(n3651), .Z(
        n1697) );
  CANR2XL U6489 ( .A(N2210), .B(n3588), .C(n3623), .D(N8145), .Z(n1702) );
  CND2XL U6490 ( .A(N5292), .B(n3695), .Z(n1701) );
  CANR2XL U6491 ( .A(mem_data1[134]), .B(n3898), .C(N8414), .D(n3651), .Z(
        n1700) );
  CANR2XL U6492 ( .A(N2209), .B(n3588), .C(n3623), .D(N8146), .Z(n1705) );
  CND2XL U6493 ( .A(N5291), .B(n3697), .Z(n1704) );
  CANR2XL U6494 ( .A(mem_data1[133]), .B(n3898), .C(N8413), .D(n3647), .Z(
        n1703) );
  CANR2XL U6495 ( .A(N2208), .B(n3588), .C(n3623), .D(N8147), .Z(n1708) );
  CND2XL U6496 ( .A(N5290), .B(n3697), .Z(n1707) );
  CANR2XL U6497 ( .A(mem_data1[132]), .B(n3898), .C(N8412), .D(n3647), .Z(
        n1706) );
  CANR2XL U6498 ( .A(N2207), .B(n3588), .C(n3623), .D(N8148), .Z(n1711) );
  CND2XL U6499 ( .A(N5289), .B(n3697), .Z(n1710) );
  CANR2XL U6500 ( .A(mem_data1[131]), .B(n3898), .C(N8411), .D(n3647), .Z(
        n1709) );
  CANR2XL U6501 ( .A(N2206), .B(n3588), .C(n3623), .D(N8149), .Z(n1714) );
  CND2XL U6502 ( .A(N5288), .B(n3697), .Z(n1713) );
  CANR2XL U6503 ( .A(mem_data1[130]), .B(n3898), .C(N8410), .D(n3647), .Z(
        n1712) );
  CANR2XL U6504 ( .A(N2205), .B(n3588), .C(n3623), .D(N8150), .Z(n1717) );
  CND2XL U6505 ( .A(N5287), .B(n3697), .Z(n1716) );
  CANR2XL U6506 ( .A(mem_data1[129]), .B(n3898), .C(N8409), .D(n3647), .Z(
        n1715) );
  CND2XL U6507 ( .A(N5286), .B(n3697), .Z(n1719) );
  CANR2XL U6508 ( .A(mem_data1[128]), .B(n3898), .C(N8408), .D(n3647), .Z(
        n1718) );
  CANR2XL U6509 ( .A(mem_data1[127]), .B(n3898), .C(N8407), .D(n3647), .Z(
        n1721) );
  CND2XL U6510 ( .A(N5285), .B(n3697), .Z(n1722) );
  CANR2XL U6511 ( .A(mem_data1[126]), .B(n3898), .C(N8406), .D(n3647), .Z(
        n1724) );
  CND2XL U6512 ( .A(N5284), .B(n3697), .Z(n1725) );
  CANR2XL U6513 ( .A(mem_data1[125]), .B(n3898), .C(N8405), .D(n3647), .Z(
        n1727) );
  CND2XL U6514 ( .A(N5283), .B(n3696), .Z(n1728) );
  CANR2XL U6515 ( .A(N2200), .B(n3589), .C(n3623), .D(N8155), .Z(n1732) );
  CND2XL U6516 ( .A(N5282), .B(n3697), .Z(n1731) );
  CANR2XL U6517 ( .A(mem_data1[124]), .B(n3898), .C(N8404), .D(n3647), .Z(
        n1730) );
  CANR2XL U6518 ( .A(mem_data1[122]), .B(n3898), .C(N8402), .D(n3647), .Z(
        n1736) );
  CND2XL U6519 ( .A(N5280), .B(n3697), .Z(n1737) );
  CANR2XL U6520 ( .A(mem_data1[121]), .B(n3898), .C(N8401), .D(n3647), .Z(
        n1739) );
  CND2XL U6521 ( .A(N5279), .B(n3697), .Z(n1740) );
  CANR2XL U6522 ( .A(mem_data1[114]), .B(n3898), .C(N8394), .D(n3646), .Z(
        n1760) );
  CND2XL U6523 ( .A(N5272), .B(n3696), .Z(n1761) );
  CND2XL U6524 ( .A(N5271), .B(n3696), .Z(n1764) );
  CANR2XL U6525 ( .A(N2189), .B(n3589), .C(n3624), .D(N8166), .Z(n1765) );
  CND2XL U6526 ( .A(N5270), .B(n3696), .Z(n1767) );
  CANR2XL U6527 ( .A(N2188), .B(n3589), .C(n3624), .D(N8167), .Z(n1768) );
  CND2XL U6528 ( .A(N5269), .B(n3689), .Z(n1770) );
  CANR2XL U6529 ( .A(N2187), .B(n3589), .C(n3624), .D(N8168), .Z(n1771) );
  CANR2XL U6530 ( .A(mem_data1[109]), .B(n3898), .C(N8389), .D(n3646), .Z(
        n1775) );
  CND2XL U6531 ( .A(N5267), .B(n3683), .Z(n1776) );
  CANR2XL U6532 ( .A(N2184), .B(n3589), .C(n3624), .D(N8171), .Z(n1780) );
  CND2XL U6533 ( .A(N5266), .B(n3686), .Z(n1779) );
  CANR2XL U6534 ( .A(mem_data1[108]), .B(n3898), .C(N8388), .D(n3646), .Z(
        n1778) );
  CANR2XL U6535 ( .A(N2183), .B(n3589), .C(n3624), .D(N8172), .Z(n1783) );
  CND2XL U6536 ( .A(N5265), .B(n3683), .Z(n1782) );
  CANR2XL U6537 ( .A(mem_data1[107]), .B(n3898), .C(N8387), .D(n3646), .Z(
        n1781) );
  CANR2XL U6538 ( .A(N2182), .B(n3589), .C(n3624), .D(N8173), .Z(n1786) );
  CND2XL U6539 ( .A(N5264), .B(n3689), .Z(n1785) );
  CANR2XL U6540 ( .A(mem_data1[106]), .B(n3898), .C(N8386), .D(n3646), .Z(
        n1784) );
  CANR2XL U6541 ( .A(N2181), .B(n3589), .C(n3624), .D(N8174), .Z(n1789) );
  CND2XL U6542 ( .A(N5263), .B(n3694), .Z(n1788) );
  CANR2XL U6543 ( .A(mem_data1[105]), .B(n3898), .C(N8385), .D(n3646), .Z(
        n1787) );
  CANR2XL U6544 ( .A(mem_data1[104]), .B(n3898), .C(N8384), .D(n3646), .Z(
        n1790) );
  CND2XL U6545 ( .A(N5262), .B(n3684), .Z(n1791) );
  CANR2XL U6546 ( .A(mem_data1[103]), .B(n3898), .C(N8383), .D(n3646), .Z(
        n1793) );
  CND2XL U6547 ( .A(N5261), .B(n3691), .Z(n1794) );
  CANR2XL U6548 ( .A(mem_data1[101]), .B(n3898), .C(N8381), .D(n3646), .Z(
        n1799) );
  CND2XL U6549 ( .A(N5259), .B(n3697), .Z(n1800) );
  CANR2XL U6550 ( .A(N2176), .B(n3590), .C(n3623), .D(N8179), .Z(n1804) );
  CND2XL U6551 ( .A(N5258), .B(n3689), .Z(n1803) );
  CANR2XL U6552 ( .A(mem_data1[100]), .B(n3898), .C(N8380), .D(n3646), .Z(
        n1802) );
  CANR2XL U6553 ( .A(mem_data1[99]), .B(n3898), .C(N8379), .D(n3646), .Z(n1805) );
  CND2XL U6554 ( .A(N5257), .B(n3691), .Z(n1806) );
  CND2XL U6555 ( .A(N5256), .B(n3684), .Z(n1809) );
  CANR2XL U6556 ( .A(N2174), .B(n3590), .C(n3623), .D(N8181), .Z(n1810) );
  CANR2XL U6557 ( .A(mem_data1[97]), .B(n3898), .C(N8377), .D(n3646), .Z(n1811) );
  CND2XL U6558 ( .A(N5255), .B(n3685), .Z(n1812) );
  CND2XL U6559 ( .A(N5254), .B(n3697), .Z(n1815) );
  CANR2XL U6560 ( .A(mem_data1[96]), .B(n3898), .C(N8376), .D(n3646), .Z(n1814) );
  CANR2XL U6561 ( .A(N2171), .B(n3590), .C(n3623), .D(N8184), .Z(n1819) );
  CND2XL U6562 ( .A(N5253), .B(n3697), .Z(n1818) );
  CANR2XL U6563 ( .A(mem_data1[95]), .B(n3898), .C(N8375), .D(n3646), .Z(n1817) );
  CANR2XL U6564 ( .A(N2169), .B(n3590), .C(n3623), .D(N8186), .Z(n1825) );
  CND2XL U6565 ( .A(N5251), .B(n3697), .Z(n1824) );
  CANR2XL U6566 ( .A(mem_data1[93]), .B(n3898), .C(N8373), .D(n3646), .Z(n1823) );
  CANR2XL U6567 ( .A(N2168), .B(n3590), .C(n3623), .D(N8187), .Z(n1828) );
  CND2XL U6568 ( .A(N5250), .B(n3697), .Z(n1827) );
  CANR2XL U6569 ( .A(mem_data1[92]), .B(n3898), .C(N8372), .D(n3646), .Z(n1826) );
  CANR2XL U6570 ( .A(N2167), .B(n3590), .C(n3623), .D(N8188), .Z(n1831) );
  CND2XL U6571 ( .A(N5249), .B(n3697), .Z(n1830) );
  CANR2XL U6572 ( .A(mem_data1[91]), .B(n3898), .C(N8371), .D(n3646), .Z(n1829) );
  CND2XL U6573 ( .A(N5248), .B(n3697), .Z(n1833) );
  CANR2XL U6574 ( .A(N2166), .B(n3590), .C(n3623), .D(N8189), .Z(n1834) );
  CANR2XL U6575 ( .A(N2164), .B(n3590), .C(n3625), .D(N8191), .Z(n1840) );
  CND2XL U6576 ( .A(N5246), .B(n3690), .Z(n1839) );
  CANR2XL U6577 ( .A(mem_data1[88]), .B(n3898), .C(N8368), .D(n3645), .Z(n1838) );
  CANR2XL U6578 ( .A(N2163), .B(n3590), .C(n3625), .D(N8192), .Z(n1843) );
  CND2XL U6579 ( .A(N5245), .B(n3685), .Z(n1842) );
  CANR2XL U6580 ( .A(mem_data1[87]), .B(n3898), .C(N8367), .D(n3645), .Z(n1841) );
  CANR2XL U6581 ( .A(N2162), .B(n3590), .C(n3625), .D(N8193), .Z(n1846) );
  CND2XL U6582 ( .A(N5244), .B(n3690), .Z(n1845) );
  CANR2XL U6583 ( .A(mem_data1[86]), .B(n3898), .C(N8366), .D(n3645), .Z(n1844) );
  CANR2XL U6584 ( .A(N2161), .B(n3589), .C(n3625), .D(N8194), .Z(n1849) );
  CND2XL U6585 ( .A(N5243), .B(n3697), .Z(n1848) );
  CANR2XL U6586 ( .A(mem_data1[85]), .B(n3898), .C(N8365), .D(n3645), .Z(n1847) );
  CANR2XL U6587 ( .A(N2160), .B(n3589), .C(n3625), .D(N8195), .Z(n1852) );
  CND2XL U6588 ( .A(N5242), .B(n3685), .Z(n1851) );
  CANR2XL U6589 ( .A(mem_data1[84]), .B(n3898), .C(N8364), .D(n3645), .Z(n1850) );
  CANR2XL U6590 ( .A(N2159), .B(n3589), .C(n3625), .D(N8196), .Z(n1855) );
  CND2XL U6591 ( .A(N5241), .B(n3690), .Z(n1854) );
  CANR2XL U6592 ( .A(mem_data1[83]), .B(n3898), .C(N8363), .D(n3645), .Z(n1853) );
  CANR2XL U6593 ( .A(N2158), .B(n3589), .C(n3624), .D(N8197), .Z(n1858) );
  CND2XL U6594 ( .A(N5240), .B(n3690), .Z(n1857) );
  CANR2XL U6595 ( .A(mem_data1[82]), .B(n3898), .C(N8362), .D(n3645), .Z(n1856) );
  CANR2XL U6596 ( .A(N2157), .B(n3589), .C(n3624), .D(N8198), .Z(n1861) );
  CND2XL U6597 ( .A(N5239), .B(n3690), .Z(n1860) );
  CANR2XL U6598 ( .A(mem_data1[81]), .B(n3898), .C(N8361), .D(n3645), .Z(n1859) );
  CANR2XL U6599 ( .A(N2156), .B(n3589), .C(n3624), .D(N8199), .Z(n1864) );
  CND2XL U6600 ( .A(N5238), .B(n3692), .Z(n1863) );
  CANR2XL U6601 ( .A(mem_data1[80]), .B(n3898), .C(N8360), .D(n3645), .Z(n1862) );
  CANR2XL U6602 ( .A(N2155), .B(n3589), .C(n3624), .D(N8200), .Z(n1867) );
  CND2XL U6603 ( .A(N5237), .B(n3698), .Z(n1866) );
  CANR2XL U6604 ( .A(mem_data1[79]), .B(n3898), .C(N8359), .D(n3645), .Z(n1865) );
  CANR2XL U6605 ( .A(N2154), .B(n3589), .C(n3624), .D(N8201), .Z(n1870) );
  CND2XL U6606 ( .A(N5236), .B(n3689), .Z(n1869) );
  CANR2XL U6607 ( .A(mem_data1[78]), .B(n3898), .C(N8358), .D(n3645), .Z(n1868) );
  CANR2XL U6608 ( .A(N2153), .B(n3589), .C(n3624), .D(N8202), .Z(n1873) );
  CND2XL U6609 ( .A(N5235), .B(n3698), .Z(n1872) );
  CANR2XL U6610 ( .A(mem_data1[77]), .B(n3898), .C(N8357), .D(n3645), .Z(n1871) );
  CANR2XL U6611 ( .A(N2152), .B(n3591), .C(n3624), .D(N8203), .Z(n1876) );
  CND2XL U6612 ( .A(N5234), .B(n3698), .Z(n1875) );
  CANR2XL U6613 ( .A(mem_data1[76]), .B(n3898), .C(N8356), .D(n3645), .Z(n1874) );
  CANR2XL U6614 ( .A(N2151), .B(n3591), .C(n3624), .D(N8204), .Z(n1879) );
  CND2XL U6615 ( .A(N5233), .B(n3688), .Z(n1878) );
  CANR2XL U6616 ( .A(mem_data1[75]), .B(n3898), .C(N8355), .D(n3645), .Z(n1877) );
  CANR2XL U6617 ( .A(N2150), .B(n3591), .C(n3624), .D(N8205), .Z(n1882) );
  CND2XL U6618 ( .A(N5232), .B(n3698), .Z(n1881) );
  CANR2XL U6619 ( .A(mem_data1[74]), .B(n3898), .C(N8354), .D(n3645), .Z(n1880) );
  CANR2XL U6620 ( .A(N2149), .B(n3591), .C(n3624), .D(N8206), .Z(n1885) );
  CND2XL U6621 ( .A(N5231), .B(n3698), .Z(n1884) );
  CANR2XL U6622 ( .A(mem_data1[73]), .B(n3898), .C(N8353), .D(n3645), .Z(n1883) );
  CANR2XL U6623 ( .A(N2148), .B(n3591), .C(n3624), .D(N8207), .Z(n1888) );
  CND2XL U6624 ( .A(N5230), .B(n3686), .Z(n1887) );
  CANR2XL U6625 ( .A(mem_data1[72]), .B(n3898), .C(N8352), .D(n3645), .Z(n1886) );
  CANR2XL U6626 ( .A(N2147), .B(n3591), .C(n3624), .D(N8208), .Z(n1891) );
  CND2XL U6627 ( .A(N5229), .B(n3698), .Z(n1890) );
  CANR2XL U6628 ( .A(mem_data1[71]), .B(n3898), .C(N8351), .D(n3646), .Z(n1889) );
  CANR2XL U6629 ( .A(N2146), .B(n3591), .C(n3624), .D(N8209), .Z(n1894) );
  CND2XL U6630 ( .A(N5228), .B(n3698), .Z(n1893) );
  CANR2XL U6631 ( .A(mem_data1[70]), .B(n3898), .C(N8350), .D(n3646), .Z(n1892) );
  CANR2XL U6632 ( .A(N2145), .B(n3591), .C(n3624), .D(N8210), .Z(n1897) );
  CND2XL U6633 ( .A(N5227), .B(n3693), .Z(n1896) );
  CANR2XL U6634 ( .A(mem_data1[69]), .B(n3898), .C(N8349), .D(n3646), .Z(n1895) );
  CANR2XL U6635 ( .A(N2144), .B(n3591), .C(n3624), .D(N8211), .Z(n1900) );
  CND2XL U6636 ( .A(N5226), .B(n3691), .Z(n1899) );
  CANR2XL U6637 ( .A(mem_data1[68]), .B(n3898), .C(N8348), .D(n3646), .Z(n1898) );
  CANR2XL U6638 ( .A(N2143), .B(n3591), .C(n3624), .D(N8212), .Z(n1903) );
  CND2XL U6639 ( .A(N5225), .B(n3691), .Z(n1902) );
  CANR2XL U6640 ( .A(mem_data1[67]), .B(n3898), .C(N8347), .D(n3644), .Z(n1901) );
  CANR2XL U6641 ( .A(N2142), .B(n3590), .C(n3624), .D(N8213), .Z(n1906) );
  CND2XL U6642 ( .A(N5224), .B(n3691), .Z(n1905) );
  CANR2XL U6643 ( .A(mem_data1[66]), .B(n3898), .C(N8346), .D(n3645), .Z(n1904) );
  CANR2XL U6644 ( .A(N2141), .B(n3590), .C(n3624), .D(N8214), .Z(n1909) );
  CND2XL U6645 ( .A(N5223), .B(n3691), .Z(n1908) );
  CANR2XL U6646 ( .A(mem_data1[65]), .B(n3898), .C(N8345), .D(n3645), .Z(n1907) );
  CND2XL U6647 ( .A(N5222), .B(n3691), .Z(n1911) );
  CANR2XL U6648 ( .A(mem_data1[64]), .B(n3898), .C(N8344), .D(n3645), .Z(n1910) );
  CANR2XL U6649 ( .A(mem_data1[63]), .B(n3898), .C(N8343), .D(n3645), .Z(n1913) );
  CND2XL U6650 ( .A(N5221), .B(n3691), .Z(n1914) );
  CANR2XL U6651 ( .A(N2138), .B(n3590), .C(n3626), .D(N8217), .Z(n1918) );
  CND2XL U6652 ( .A(N5220), .B(n3691), .Z(n1917) );
  CANR2XL U6653 ( .A(mem_data1[62]), .B(n3898), .C(n3644), .D(N8342), .Z(n1916) );
  CANR2XL U6654 ( .A(mem_data1[60]), .B(n3898), .C(n3644), .D(N8340), .Z(n1922) );
  CND2XL U6655 ( .A(N5218), .B(n3690), .Z(n1923) );
  CND2XL U6656 ( .A(N5217), .B(n3690), .Z(n1926) );
  CANR2XL U6657 ( .A(N2135), .B(n3590), .C(n3626), .D(N8220), .Z(n1927) );
  CND2XL U6658 ( .A(N5216), .B(n3685), .Z(n1929) );
  CANR2XL U6659 ( .A(N2134), .B(n3590), .C(n3626), .D(N8221), .Z(n1930) );
  CANR2XL U6660 ( .A(N2133), .B(n3590), .C(n3626), .D(N8222), .Z(n1933) );
  CND2XL U6661 ( .A(N5215), .B(n3697), .Z(n1932) );
  CANR2XL U6662 ( .A(mem_data1[57]), .B(n3898), .C(n3644), .D(N8337), .Z(n1931) );
  CANR2XL U6663 ( .A(N2132), .B(n3590), .C(n3625), .D(N8223), .Z(n1936) );
  CND2XL U6664 ( .A(N5214), .B(n3696), .Z(n1935) );
  CANR2XL U6665 ( .A(mem_data1[56]), .B(n3898), .C(n3644), .D(N8336), .Z(n1934) );
  CANR2XL U6666 ( .A(N2131), .B(n3590), .C(n3625), .D(N8224), .Z(n1939) );
  CND2XL U6667 ( .A(N5213), .B(n3685), .Z(n1938) );
  CANR2XL U6668 ( .A(mem_data1[55]), .B(n3898), .C(n3644), .D(N8335), .Z(n1937) );
  CANR2XL U6669 ( .A(N2130), .B(n3590), .C(n3625), .D(N8225), .Z(n1942) );
  CND2XL U6670 ( .A(N5212), .B(n3687), .Z(n1941) );
  CANR2XL U6671 ( .A(mem_data1[54]), .B(n3898), .C(n3644), .D(N8334), .Z(n1940) );
  CANR2XL U6672 ( .A(N2129), .B(n3590), .C(n3625), .D(N8226), .Z(n1945) );
  CND2XL U6673 ( .A(N5211), .B(n3694), .Z(n1944) );
  CANR2XL U6674 ( .A(mem_data1[53]), .B(n3898), .C(n3644), .D(N8333), .Z(n1943) );
  CANR2XL U6675 ( .A(N2128), .B(n3590), .C(n3625), .D(N8227), .Z(n1948) );
  CND2XL U6676 ( .A(N5210), .B(n3685), .Z(n1947) );
  CANR2XL U6677 ( .A(mem_data1[52]), .B(n3898), .C(n3644), .D(N8332), .Z(n1946) );
  CANR2XL U6678 ( .A(N2127), .B(n3602), .C(n3625), .D(N8228), .Z(n1951) );
  CND2XL U6679 ( .A(N5209), .B(n3697), .Z(n1950) );
  CANR2XL U6680 ( .A(mem_data1[51]), .B(n3898), .C(n3644), .D(N8331), .Z(n1949) );
  CANR2XL U6681 ( .A(N2126), .B(n3592), .C(n3625), .D(N8229), .Z(n1954) );
  CND2XL U6682 ( .A(N5208), .B(n3695), .Z(n1953) );
  CANR2XL U6683 ( .A(mem_data1[50]), .B(n3898), .C(n3644), .D(N8330), .Z(n1952) );
  CANR2XL U6684 ( .A(N2125), .B(n3592), .C(n3625), .D(N8230), .Z(n1957) );
  CND2XL U6685 ( .A(N5207), .B(n3685), .Z(n1956) );
  CANR2XL U6686 ( .A(mem_data1[49]), .B(n3898), .C(n3644), .D(N8329), .Z(n1955) );
  CANR2XL U6687 ( .A(N2124), .B(n3592), .C(n3625), .D(N8231), .Z(n1960) );
  CND2XL U6688 ( .A(N5206), .B(n3695), .Z(n1959) );
  CANR2XL U6689 ( .A(mem_data1[48]), .B(n3898), .C(n3644), .D(N8328), .Z(n1958) );
  CANR2XL U6690 ( .A(N2123), .B(n3592), .C(n3625), .D(N8232), .Z(n1963) );
  CND2XL U6691 ( .A(N5205), .B(n3690), .Z(n1962) );
  CANR2XL U6692 ( .A(mem_data1[47]), .B(n3898), .C(n3644), .D(N8327), .Z(n1961) );
  CANR2XL U6693 ( .A(mem_data1[46]), .B(n3898), .C(n3644), .D(N8326), .Z(n1964) );
  CND2XL U6694 ( .A(N5204), .B(n3685), .Z(n1965) );
  CANR2XL U6695 ( .A(N2121), .B(n3592), .C(n3625), .D(N8234), .Z(n1969) );
  CND2XL U6696 ( .A(N5203), .B(n3692), .Z(n1968) );
  CANR2XL U6697 ( .A(mem_data1[45]), .B(n3898), .C(n3644), .D(N8325), .Z(n1967) );
  CANR2XL U6698 ( .A(N2120), .B(n3592), .C(n3625), .D(N8235), .Z(n1972) );
  CND2XL U6699 ( .A(N5202), .B(n3692), .Z(n1971) );
  CANR2XL U6700 ( .A(mem_data1[44]), .B(n3898), .C(N8324), .D(n3677), .Z(n1970) );
  CANR2XL U6701 ( .A(N2119), .B(n3592), .C(n3625), .D(N8236), .Z(n1975) );
  CND2XL U6702 ( .A(N5201), .B(n3692), .Z(n1974) );
  CANR2XL U6703 ( .A(mem_data1[43]), .B(n3898), .C(N8323), .D(n3677), .Z(n1973) );
  CANR2XL U6704 ( .A(N2118), .B(n3591), .C(n3625), .D(N8237), .Z(n1978) );
  CND2XL U6705 ( .A(N5200), .B(n3692), .Z(n1977) );
  CANR2XL U6706 ( .A(mem_data1[42]), .B(n3898), .C(N8322), .D(n3677), .Z(n1976) );
  CANR2XL U6707 ( .A(N2117), .B(n3591), .C(n3625), .D(N8238), .Z(n1981) );
  CND2XL U6708 ( .A(N5199), .B(n3692), .Z(n1980) );
  CANR2XL U6709 ( .A(mem_data1[41]), .B(n3898), .C(N8321), .D(n3677), .Z(n1979) );
  CANR2XL U6710 ( .A(N2116), .B(n3591), .C(n3625), .D(N8239), .Z(n1984) );
  CND2XL U6711 ( .A(N5198), .B(n3692), .Z(n1983) );
  CANR2XL U6712 ( .A(mem_data1[40]), .B(n3898), .C(N8320), .D(n3677), .Z(n1982) );
  CANR2XL U6713 ( .A(N2115), .B(n3591), .C(n3625), .D(N8240), .Z(n1987) );
  CND2XL U6714 ( .A(N5197), .B(n3691), .Z(n1986) );
  CANR2XL U6715 ( .A(mem_data1[39]), .B(n3898), .C(N8319), .D(n3676), .Z(n1985) );
  CANR2XL U6716 ( .A(N2114), .B(n3591), .C(n3625), .D(N8241), .Z(n1990) );
  CND2XL U6717 ( .A(N5196), .B(n3691), .Z(n1989) );
  CANR2XL U6718 ( .A(mem_data1[38]), .B(n3898), .C(N8318), .D(n3677), .Z(n1988) );
  CANR2XL U6719 ( .A(N2113), .B(n3591), .C(n3625), .D(N8242), .Z(n1993) );
  CND2XL U6720 ( .A(N5195), .B(n3691), .Z(n1992) );
  CANR2XL U6721 ( .A(mem_data1[37]), .B(n3898), .C(N8317), .D(n3677), .Z(n1991) );
  CANR2XL U6722 ( .A(N2112), .B(n3591), .C(n3625), .D(N8243), .Z(n1996) );
  CND2XL U6723 ( .A(N5194), .B(n3691), .Z(n1995) );
  CANR2XL U6724 ( .A(mem_data1[36]), .B(n3898), .C(N8316), .D(n3677), .Z(n1994) );
  CANR2XL U6725 ( .A(mem_data1[35]), .B(n3898), .C(N8315), .D(n3677), .Z(n1997) );
  CND2XL U6726 ( .A(N5193), .B(n3691), .Z(n1998) );
  CANR2XL U6727 ( .A(N2110), .B(n3591), .C(n3636), .D(N8245), .Z(n2002) );
  CND2XL U6728 ( .A(N5192), .B(n3691), .Z(n2001) );
  CANR2XL U6729 ( .A(mem_data1[34]), .B(n3898), .C(N8314), .D(n3677), .Z(n2000) );
  CND2XL U6730 ( .A(N5191), .B(n3691), .Z(n2004) );
  CANR2XL U6731 ( .A(N2109), .B(n3591), .C(n3635), .D(N8246), .Z(n2005) );
  CANR2XL U6732 ( .A(N2108), .B(n3591), .C(n3636), .D(N8247), .Z(n2008) );
  CND2XL U6733 ( .A(N5190), .B(n3691), .Z(n2007) );
  CANR2XL U6734 ( .A(mem_data1[32]), .B(n3898), .C(N8312), .D(n3677), .Z(n2006) );
  CANR2XL U6735 ( .A(N2107), .B(n3591), .C(n3636), .D(N8248), .Z(n2011) );
  CND2XL U6736 ( .A(N5189), .B(n3691), .Z(n2010) );
  CANR2XL U6737 ( .A(mem_data1[31]), .B(n3898), .C(N8311), .D(n3677), .Z(n2009) );
  CANR2XL U6738 ( .A(N2106), .B(n3591), .C(n3623), .D(N8249), .Z(n2014) );
  CND2XL U6739 ( .A(N5188), .B(n3691), .Z(n2013) );
  CANR2XL U6740 ( .A(mem_data1[30]), .B(n3898), .C(N8310), .D(n3677), .Z(n2012) );
  CANR2XL U6741 ( .A(N2105), .B(n3590), .C(n3627), .D(N8250), .Z(n2017) );
  CND2XL U6742 ( .A(N5187), .B(n3691), .Z(n2016) );
  CANR2XL U6743 ( .A(mem_data1[29]), .B(n3898), .C(N8309), .D(n3677), .Z(n2015) );
  CANR2XL U6744 ( .A(N2104), .B(n3592), .C(n3627), .D(N8251), .Z(n2020) );
  CND2XL U6745 ( .A(N5186), .B(n3691), .Z(n2019) );
  CANR2XL U6746 ( .A(mem_data1[28]), .B(n3898), .C(N8308), .D(n3677), .Z(n2018) );
  CANR2XL U6747 ( .A(N2103), .B(n3592), .C(n3627), .D(N8252), .Z(n2023) );
  CND2XL U6748 ( .A(N5185), .B(n3691), .Z(n2022) );
  CANR2XL U6749 ( .A(mem_data1[27]), .B(n3898), .C(N8307), .D(n3677), .Z(n2021) );
  CANR2XL U6750 ( .A(N2102), .B(n3592), .C(n3627), .D(N8253), .Z(n2026) );
  CND2XL U6751 ( .A(N5184), .B(n3691), .Z(n2025) );
  CANR2XL U6752 ( .A(mem_data1[26]), .B(n3898), .C(N8306), .D(n3677), .Z(n2024) );
  CANR2XL U6753 ( .A(N2101), .B(n3592), .C(n3627), .D(N8254), .Z(n2029) );
  CND2XL U6754 ( .A(N5183), .B(n3691), .Z(n2028) );
  CANR2XL U6755 ( .A(mem_data1[25]), .B(n3898), .C(N8305), .D(n3677), .Z(n2027) );
  CANR2XL U6756 ( .A(N2100), .B(n3592), .C(n3627), .D(N8255), .Z(n2032) );
  CND2XL U6757 ( .A(N5182), .B(n3691), .Z(n2031) );
  CANR2XL U6758 ( .A(mem_data1[24]), .B(n3898), .C(N8304), .D(n3675), .Z(n2030) );
  CANR2XL U6759 ( .A(N2099), .B(n3592), .C(n3627), .D(N8256), .Z(n2035) );
  CND2XL U6760 ( .A(N5181), .B(n3686), .Z(n2034) );
  CANR2XL U6761 ( .A(mem_data1[23]), .B(n3898), .C(N8303), .D(n3675), .Z(n2033) );
  CANR2XL U6762 ( .A(N2098), .B(n3592), .C(n3627), .D(N8257), .Z(n2038) );
  CND2XL U6763 ( .A(N5180), .B(n3691), .Z(n2037) );
  CANR2XL U6764 ( .A(mem_data1[22]), .B(n3898), .C(N8302), .D(n3675), .Z(n2036) );
  CANR2XL U6765 ( .A(N2097), .B(n3592), .C(n3627), .D(N8258), .Z(n2041) );
  CND2XL U6766 ( .A(N5179), .B(n3687), .Z(n2040) );
  CANR2XL U6767 ( .A(mem_data1[21]), .B(n3898), .C(N8301), .D(n3675), .Z(n2039) );
  CANR2XL U6768 ( .A(N2096), .B(n3594), .C(n3627), .D(N8259), .Z(n2044) );
  CND2XL U6769 ( .A(N5178), .B(n3691), .Z(n2043) );
  CANR2XL U6770 ( .A(mem_data1[20]), .B(n3898), .C(N8300), .D(n3675), .Z(n2042) );
  CANR2XL U6771 ( .A(N2095), .B(n3596), .C(n3626), .D(N8260), .Z(n2047) );
  CND2XL U6772 ( .A(N5177), .B(n3693), .Z(n2046) );
  CANR2XL U6773 ( .A(mem_data1[19]), .B(n3898), .C(N8299), .D(n3675), .Z(n2045) );
  CANR2XL U6774 ( .A(N2094), .B(n3570), .C(n3627), .D(N8261), .Z(n2050) );
  CND2XL U6775 ( .A(N5176), .B(n3691), .Z(n2049) );
  CANR2XL U6776 ( .A(mem_data1[18]), .B(n3898), .C(N8298), .D(n3675), .Z(n2048) );
  CANR2XL U6777 ( .A(N2093), .B(n3593), .C(n3626), .D(N8262), .Z(n2053) );
  CND2XL U6778 ( .A(N5175), .B(n3694), .Z(n2052) );
  CANR2XL U6779 ( .A(mem_data1[17]), .B(n3898), .C(N8297), .D(n3676), .Z(n2051) );
  CANR2XL U6780 ( .A(N2092), .B(n3593), .C(n3626), .D(N8263), .Z(n2056) );
  CND2XL U6781 ( .A(N5174), .B(n3692), .Z(n2055) );
  CANR2XL U6782 ( .A(mem_data1[16]), .B(n3898), .C(N8296), .D(n3676), .Z(n2054) );
  CANR2XL U6783 ( .A(N2091), .B(n3593), .C(n3626), .D(N8264), .Z(n2059) );
  CND2XL U6784 ( .A(N5173), .B(n3692), .Z(n2058) );
  CANR2XL U6785 ( .A(mem_data1[15]), .B(n3898), .C(N8295), .D(n3676), .Z(n2057) );
  CANR2XL U6786 ( .A(N2752), .B(n3583), .C(n3618), .D(N7603), .Z(n3169) );
  CND2XL U6787 ( .A(N5834), .B(n3691), .Z(n3168) );
  CANR2XL U6788 ( .A(mem_data1[676]), .B(n3898), .C(N8956), .D(n3665), .Z(
        n3167) );
  CANR2XL U6789 ( .A(n3898), .B(mem_data1[14]), .C(N8294), .D(n3676), .Z(n2060) );
  CND2XL U6790 ( .A(N5172), .B(n3692), .Z(n2061) );
  CANR2XL U6791 ( .A(N2089), .B(n3593), .C(n3626), .D(N8266), .Z(n2065) );
  CND2XL U6792 ( .A(N5171), .B(n3692), .Z(n2064) );
  CANR2XL U6793 ( .A(n3898), .B(mem_data1[13]), .C(N8293), .D(n3676), .Z(n2063) );
  CANR2XL U6794 ( .A(N2088), .B(n3593), .C(n3627), .D(N8267), .Z(n2068) );
  CND2XL U6795 ( .A(N5170), .B(n3692), .Z(n2067) );
  CANR2XL U6796 ( .A(n3898), .B(mem_data1[12]), .C(N8292), .D(n3675), .Z(n2066) );
  CANR2XL U6797 ( .A(N2087), .B(n3593), .C(n3626), .D(N8268), .Z(n2071) );
  CND2XL U6798 ( .A(N5169), .B(n3692), .Z(n2070) );
  CANR2XL U6799 ( .A(n3898), .B(mem_data1[11]), .C(N8291), .D(n3676), .Z(n2069) );
  CANR2XL U6800 ( .A(N2086), .B(n3593), .C(n3626), .D(N8269), .Z(n2074) );
  CND2XL U6801 ( .A(N5168), .B(n3692), .Z(n2073) );
  CANR2XL U6802 ( .A(n3898), .B(mem_data1[10]), .C(N8290), .D(n3676), .Z(n2072) );
  CANR2XL U6803 ( .A(N2085), .B(n3593), .C(n3628), .D(N8270), .Z(n2077) );
  CND2XL U6804 ( .A(N5167), .B(n3692), .Z(n2076) );
  CANR2XL U6805 ( .A(n3898), .B(mem_data1[9]), .C(N8289), .D(n3676), .Z(n2075)
         );
  CANR2XL U6806 ( .A(N2084), .B(n3593), .C(n3626), .D(N8271), .Z(n2080) );
  CND2XL U6807 ( .A(N5166), .B(n3692), .Z(n2079) );
  CANR2XL U6808 ( .A(n3898), .B(mem_data1[8]), .C(N8288), .D(n3676), .Z(n2078)
         );
  CANR2XL U6809 ( .A(N2083), .B(n3593), .C(n3626), .D(N8272), .Z(n2083) );
  CND2XL U6810 ( .A(N5165), .B(n3692), .Z(n2082) );
  CANR2XL U6811 ( .A(n3898), .B(mem_data1[7]), .C(N8287), .D(n3676), .Z(n2081)
         );
  CND2XL U6812 ( .A(N5164), .B(n3692), .Z(n2085) );
  CANR2XL U6813 ( .A(n3898), .B(mem_data1[6]), .C(N8286), .D(n3676), .Z(n2084)
         );
  CND2XL U6814 ( .A(N5163), .B(n3692), .Z(n2088) );
  CANR2XL U6815 ( .A(n3898), .B(mem_data1[5]), .C(N8285), .D(n3676), .Z(n2087)
         );
  CND2XL U6816 ( .A(N5162), .B(n3692), .Z(n2091) );
  CANR2XL U6817 ( .A(N2080), .B(n3593), .C(n3628), .D(N8275), .Z(n2092) );
  CND2XL U6818 ( .A(N5161), .B(n3692), .Z(n2094) );
  CANR2XL U6819 ( .A(n3898), .B(mem_data1[3]), .C(N8283), .D(n3677), .Z(n2093)
         );
  CND2XL U6820 ( .A(N5160), .B(n3692), .Z(n2097) );
  CANR2XL U6821 ( .A(n3898), .B(mem_data1[2]), .C(N8282), .D(n3677), .Z(n2096)
         );
  CND2XL U6822 ( .A(N5159), .B(n3693), .Z(n2100) );
  CANR2XL U6823 ( .A(n3898), .B(mem_data1[1]), .C(N8281), .D(n3674), .Z(n2099)
         );
  CND2XL U6824 ( .A(N5158), .B(n3693), .Z(n2103) );
  CANR2XL U6825 ( .A(n3898), .B(mem_data1[0]), .C(N8280), .D(n3674), .Z(n2102)
         );
  CANR2XL U6826 ( .A(n3698), .B(N8266), .C(mem_data1[13]), .D(n3250), .Z(n59)
         );
  CANR2XL U6827 ( .A(n3698), .B(N8267), .C(mem_data1[12]), .D(n3250), .Z(n60)
         );
  CANR2XL U6828 ( .A(n3698), .B(N8268), .C(mem_data1[11]), .D(n3250), .Z(n61)
         );
  CANR2XL U6829 ( .A(n3698), .B(N8269), .C(mem_data1[10]), .D(n3250), .Z(n62)
         );
  CANR2XL U6830 ( .A(n3698), .B(N8270), .C(mem_data1[9]), .D(n3250), .Z(n63)
         );
  CANR2XL U6831 ( .A(n3698), .B(N8271), .C(mem_data1[8]), .D(n3250), .Z(n64)
         );
  CANR2XL U6832 ( .A(n3698), .B(N8272), .C(mem_data1[7]), .D(n3250), .Z(n65)
         );
  CANR2XL U6833 ( .A(n3698), .B(N8273), .C(mem_data1[6]), .D(n3250), .Z(n66)
         );
  CANR2XL U6834 ( .A(n3698), .B(N8274), .C(mem_data1[5]), .D(n3250), .Z(n67)
         );
  CANR2XL U6835 ( .A(n3698), .B(N8275), .C(mem_data1[4]), .D(n3250), .Z(n68)
         );
  CANR2XL U6836 ( .A(n3698), .B(N8276), .C(mem_data1[3]), .D(n3250), .Z(n69)
         );
  CANR2XL U6837 ( .A(n3698), .B(N8277), .C(mem_data1[2]), .D(n3250), .Z(n70)
         );
  CANR2XL U6838 ( .A(n3698), .B(N8278), .C(mem_data1[1]), .D(n3250), .Z(n71)
         );
  CANR2XL U6839 ( .A(n3698), .B(N8279), .C(mem_data1[0]), .D(n3250), .Z(n72)
         );
  CANR2XL U6840 ( .A(N6222), .B(n2105), .C(N2066), .D(n3898), .Z(n2125) );
  CND2XL U6841 ( .A(n2124), .B(n2125), .Z(N10348) );
  CNIVX4 U6842 ( .A(lenin0[3]), .Z(n3897) );
  CNIVX4 U6843 ( .A(N2068), .Z(n3896) );
  CNR2XL U6844 ( .A(n3834), .B(n5844), .Z(N23) );
  CNR2XL U6845 ( .A(n3836), .B(n5374), .Z(N21) );
  CNR2XL U6846 ( .A(n3851), .B(n6225), .Z(N25) );
  CNIVXL U6847 ( .A(N2069), .Z(n3753) );
  CENX1 U6848 ( .A(n3251), .B(mem_data1[132]), .Z(N8147) );
  COR2X1 U6849 ( .A(n3829), .B(n5568), .Z(n3251) );
  CNR2XL U6850 ( .A(n3818), .B(n4767), .Z(N159) );
  CNR2XL U6851 ( .A(n3822), .B(n4766), .Z(N158) );
  CNR2XL U6852 ( .A(n3832), .B(n4763), .Z(N157) );
  CNR2XL U6853 ( .A(n3816), .B(n6515), .Z(N155) );
  CND2XL U6854 ( .A(n4856), .B(n3726), .Z(n4709) );
  CND2XL U6855 ( .A(n4852), .B(n3727), .Z(n4699) );
  CND2XL U6856 ( .A(n4850), .B(n3724), .Z(n4695) );
  CND2XL U6857 ( .A(n4848), .B(n3728), .Z(n4691) );
  CND2XL U6858 ( .A(n4833), .B(n3728), .Z(n4653) );
  CND2XL U6859 ( .A(n4843), .B(n3724), .Z(n4682) );
  CEOX1 U6860 ( .A(n3252), .B(mem_data1[446]), .Z(N7833) );
  CND2XL U6861 ( .A(n4871), .B(n3726), .Z(n4737) );
  CND2XL U6862 ( .A(n4869), .B(n3725), .Z(n4733) );
  CND2XL U6863 ( .A(n4866), .B(n3724), .Z(n4729) );
  CND2XL U6864 ( .A(n4845), .B(n3729), .Z(n4688) );
  CEOX1 U6865 ( .A(n3253), .B(mem_data1[417]), .Z(N7862) );
  CNR2X1 U6866 ( .A(n3821), .B(n5393), .Z(n3253) );
  CEOX1 U6867 ( .A(n3254), .B(mem_data1[444]), .Z(N7835) );
  CEOX1 U6868 ( .A(n3255), .B(mem_data1[443]), .Z(N7836) );
  CEOX1 U6869 ( .A(n3256), .B(mem_data1[442]), .Z(N7837) );
  CEOX1 U6870 ( .A(n3257), .B(mem_data1[441]), .Z(N7838) );
  CEOX1 U6871 ( .A(n3258), .B(mem_data1[437]), .Z(N7842) );
  CEOX1 U6872 ( .A(n3259), .B(mem_data1[436]), .Z(N7843) );
  CEOX1 U6873 ( .A(n3260), .B(mem_data1[419]), .Z(N7860) );
  CNR2X1 U6874 ( .A(n3825), .B(n5395), .Z(n3260) );
  CEOX1 U6875 ( .A(n3261), .B(mem_data1[300]), .Z(N7979) );
  CNR2X1 U6876 ( .A(n3853), .B(n5405), .Z(n3261) );
  CEOX1 U6877 ( .A(n3262), .B(mem_data1[298]), .Z(N7981) );
  CNR2X1 U6878 ( .A(n5403), .B(n3850), .Z(n3262) );
  CEOX1 U6879 ( .A(n3263), .B(mem_data1[291]), .Z(N7988) );
  CNR2X1 U6880 ( .A(n3848), .B(n5395), .Z(n3263) );
  CND2XL U6881 ( .A(n4841), .B(n3728), .Z(n4676) );
  CND2XL U6882 ( .A(n4862), .B(n3724), .Z(n4721) );
  CND2XL U6883 ( .A(n4864), .B(n3729), .Z(n4725) );
  CND2XL U6884 ( .A(n4858), .B(n3725), .Z(n4713) );
  CND2XL U6885 ( .A(n4854), .B(n3721), .Z(n4703) );
  CND2XL U6886 ( .A(n4839), .B(n3730), .Z(n4670) );
  CND2XL U6887 ( .A(n4837), .B(n3726), .Z(n4667) );
  CND2XL U6888 ( .A(n4831), .B(n3727), .Z(n4647) );
  CND2XL U6889 ( .A(n4829), .B(n3729), .Z(n4641) );
  CND2XL U6890 ( .A(n4824), .B(n3723), .Z(n4621) );
  CNR2XL U6891 ( .A(n5096), .B(N2066), .Z(n5107) );
  CNR2XL U6892 ( .A(n5660), .B(N2066), .Z(n5671) );
  CNR2XL U6893 ( .A(n4535), .B(N2066), .Z(n4589) );
  CNR2XL U6894 ( .A(n4441), .B(N2066), .Z(n4475) );
  CNR2IXL U6895 ( .B(n4756), .A(n3199), .Z(n4819) );
  CNR2IXL U6896 ( .B(n4764), .A(n3215), .Z(n4832) );
  CNR2IXL U6897 ( .B(n6206), .A(n3209), .Z(n6273) );
  CIVDXL U6898 ( .A(wr_ptr[7]), .Z0(n3813), .Z1(n3814) );
  CND2XL U6899 ( .A(n5750), .B(n3201), .Z(n5816) );
  CAN2XL U6900 ( .A(datain0[30]), .B(n4389), .Z(n5647) );
  CAN2XL U6901 ( .A(datain0[31]), .B(n4389), .Z(n5654) );
  CAN2XL U6902 ( .A(datain0[12]), .B(n4388), .Z(n5522) );
  CAN2XL U6903 ( .A(datain0[28]), .B(n4388), .Z(n5632) );
  CAN2XL U6904 ( .A(datain0[29]), .B(n4389), .Z(n5640) );
  CEOX1 U6905 ( .A(n3264), .B(mem_data1[293]), .Z(N7986) );
  CIVDXL U6906 ( .A(lenin0[2]), .Z0(n3769), .Z1(n3770) );
  COR2X1 U6907 ( .A(n3898), .B(N10358), .Z(n55) );
  CMXI2X1 U6908 ( .A0(n15076), .A1(n4426), .S(n3804), .Z(n15078) );
  CMXI2X1 U6909 ( .A0(n14408), .A1(n4427), .S(n3804), .Z(n14410) );
  CNR2X1 U6910 ( .A(n4215), .B(n6059), .Z(n6079) );
  CNR2X1 U6911 ( .A(n4214), .B(n6054), .Z(n6075) );
  CNR2X1 U6912 ( .A(n4216), .B(n5490), .Z(n5514) );
  CNR2X1 U6913 ( .A(n4216), .B(n4933), .Z(n4957) );
  CNR2X1 U6914 ( .A(n4212), .B(n5495), .Z(n5520) );
  CNR2X1 U6915 ( .A(n4215), .B(n4640), .Z(n4687) );
  CNR2IX1 U6916 ( .B(n6223), .A(n3214), .Z(n6291) );
  CNR2IX1 U6917 ( .B(n6213), .A(n3206), .Z(n6280) );
  CNR2IX1 U6918 ( .B(n6211), .A(n3200), .Z(n6278) );
  CNR2IX1 U6919 ( .B(n6215), .A(n3200), .Z(n6282) );
  CNR2IX1 U6920 ( .B(n6221), .A(n3212), .Z(n6289) );
  CNR2IX1 U6921 ( .B(n4796), .A(n3202), .Z(n4862) );
  CNR2IX1 U6922 ( .B(n4794), .A(n3200), .Z(n4860) );
  CNR2IX1 U6923 ( .B(n6219), .A(n3206), .Z(n6286) );
  CNR2IX1 U6924 ( .B(n6209), .A(n3208), .Z(n6276) );
  CNR2IX1 U6925 ( .B(n6198), .A(n3212), .Z(n6265) );
  CNR2IX1 U6926 ( .B(n4786), .A(n3212), .Z(n4852) );
  CNR2IX1 U6927 ( .B(n4783), .A(n3212), .Z(n4850) );
  CNR2IX1 U6928 ( .B(n4781), .A(n3216), .Z(n4848) );
  CNR2IX1 U6929 ( .B(n4779), .A(n3202), .Z(n4845) );
  CNR2IX1 U6930 ( .B(n4773), .A(n3206), .Z(n4839) );
  CNR2IX1 U6931 ( .B(n6196), .A(n3212), .Z(n6263) );
  CNR2IX1 U6932 ( .B(n6202), .A(n3204), .Z(n6270) );
  CNR2IX1 U6933 ( .B(n6207), .A(n3204), .Z(n6274) );
  CNR2IX1 U6934 ( .B(n6205), .A(n3202), .Z(n6272) );
  CNR2IX1 U6935 ( .B(n6188), .A(n3214), .Z(n6255) );
  CNR2IX1 U6936 ( .B(n6190), .A(n3214), .Z(n6257) );
  CNR2IX1 U6937 ( .B(n6200), .A(n3210), .Z(n6268) );
  CNR2IX1 U6938 ( .B(n4777), .A(n3204), .Z(n4843) );
  CNR2IX1 U6939 ( .B(n4769), .A(n3204), .Z(n4835) );
  CNR2IX1 U6940 ( .B(n4743), .A(n3200), .Z(n4831) );
  CNR2IX1 U6941 ( .B(n4759), .A(n3206), .Z(n4822) );
  CNR2IX1 U6942 ( .B(n4757), .A(n3208), .Z(n4820) );
  CNR2IX1 U6943 ( .B(n4755), .A(n3210), .Z(n4818) );
  CNR2IX1 U6944 ( .B(n4753), .A(n3212), .Z(n4816) );
  CNR2IX1 U6945 ( .B(n4751), .A(n3204), .Z(n4814) );
  CNR2IX1 U6946 ( .B(n6194), .A(n3216), .Z(n6261) );
  CNR2IX1 U6947 ( .B(n6192), .A(n3210), .Z(n6259) );
  CNR2IX1 U6948 ( .B(n6186), .A(n3208), .Z(n6253) );
  CNR2IX1 U6949 ( .B(n6184), .A(n3214), .Z(n6251) );
  CNR2IX1 U6950 ( .B(n6181), .A(n3210), .Z(n6249) );
  CNR2IX1 U6951 ( .B(n6179), .A(n3216), .Z(n6247) );
  CNR2IX1 U6952 ( .B(n6177), .A(n3208), .Z(n6244) );
  CNR2IX1 U6953 ( .B(n6175), .A(n3202), .Z(n6242) );
  CNR2IX1 U6954 ( .B(n6176), .A(n3213), .Z(n6243) );
  CNR2IX1 U6955 ( .B(n6174), .A(n3209), .Z(n6241) );
  CNR2IX1 U6956 ( .B(n4654), .A(n3213), .Z(n4826) );
  CNR2IX1 U6957 ( .B(n4760), .A(n3213), .Z(n4823) );
  CNR2IX1 U6958 ( .B(n4754), .A(n3199), .Z(n4817) );
  CNR2IX1 U6959 ( .B(n4752), .A(n3203), .Z(n4815) );
  CNR2IX1 U6960 ( .B(n6191), .A(n3203), .Z(n6258) );
  CNR2IX1 U6961 ( .B(n6193), .A(n3205), .Z(n6260) );
  CNR2IX1 U6962 ( .B(n6187), .A(n3211), .Z(n6254) );
  CNR2IX1 U6963 ( .B(n4776), .A(n3209), .Z(n4842) );
  CNR2IX1 U6964 ( .B(n4768), .A(n3209), .Z(n4834) );
  CNR2IX1 U6965 ( .B(n4742), .A(n3209), .Z(n4830) );
  CNR2IX1 U6966 ( .B(n4704), .A(n3213), .Z(n4828) );
  CNR2IX1 U6967 ( .B(n4750), .A(n3199), .Z(n4813) );
  CNR2IX1 U6968 ( .B(n6197), .A(n3215), .Z(n6264) );
  CNR2IX1 U6969 ( .B(n6189), .A(n3199), .Z(n6256) );
  CNR2IX1 U6970 ( .B(n6199), .A(n3207), .Z(n6267) );
  CNR2IX1 U6971 ( .B(n6195), .A(n3211), .Z(n6262) );
  CNR2IX1 U6972 ( .B(n6204), .A(n3201), .Z(n6271) );
  CNR2IX1 U6973 ( .B(n6201), .A(n3211), .Z(n6269) );
  CNR2IX1 U6974 ( .B(n6218), .A(n3199), .Z(n6285) );
  CNR2IX1 U6975 ( .B(n6208), .A(n3205), .Z(n6275) );
  CNR2IX1 U6976 ( .B(n4789), .A(n3213), .Z(n4855) );
  CNR2IX1 U6977 ( .B(n4787), .A(n3201), .Z(n4853) );
  CNR2IX1 U6978 ( .B(n6216), .A(n3211), .Z(n6283) );
  CNR2IX1 U6979 ( .B(n4803), .A(n3209), .Z(n4870) );
  CNR2IX1 U6980 ( .B(n4801), .A(n3205), .Z(n4868) );
  CNR2IX1 U6981 ( .B(n4799), .A(n3201), .Z(n4865) );
  CNR2IX1 U6982 ( .B(n4797), .A(n3203), .Z(n4863) );
  CNR2IX1 U6983 ( .B(n4795), .A(n3201), .Z(n4861) );
  CNR2IX1 U6984 ( .B(n4793), .A(n3201), .Z(n4859) );
  CNR2IX1 U6985 ( .B(n4791), .A(n3211), .Z(n4857) );
  CNR2IX1 U6986 ( .B(n4785), .A(n3215), .Z(n4851) );
  CNR2IX1 U6987 ( .B(n4782), .A(n3215), .Z(n4849) );
  CNR2IX1 U6988 ( .B(n4780), .A(n3205), .Z(n4847) );
  CNR2IX1 U6989 ( .B(n4778), .A(n3207), .Z(n4844) );
  CNR2IX1 U6990 ( .B(n4774), .A(n3203), .Z(n4840) );
  CNR2IX1 U6991 ( .B(n4772), .A(n3213), .Z(n4838) );
  CNR2IX1 U6992 ( .B(n6220), .A(n3215), .Z(n6288) );
  CNR2IX1 U6993 ( .B(n6222), .A(n3205), .Z(n6290) );
  CNR2X1 U6994 ( .A(n3506), .B(n12719), .Z(N9302) );
  CNR2X1 U6995 ( .A(n3505), .B(n12720), .Z(N9303) );
  CNR2X1 U6996 ( .A(n3416), .B(n6574), .Z(N3097) );
  CNR2X1 U6997 ( .A(n3504), .B(n6573), .Z(N3096) );
  CNR2X1 U6998 ( .A(n3514), .B(n6572), .Z(N3095) );
  CNR2X1 U6999 ( .A(n3503), .B(n6571), .Z(N3094) );
  CNR2X1 U7000 ( .A(n3513), .B(n6570), .Z(N3093) );
  CNR2X1 U7001 ( .A(n3512), .B(n6569), .Z(N3092) );
  CNR2X1 U7002 ( .A(n3270), .B(n9647), .Z(N6180) );
  CNR2X1 U7003 ( .A(n3270), .B(n9648), .Z(N6181) );
  CNR2IX1 U7004 ( .B(n4792), .A(n3202), .Z(n4858) );
  CNR2IX1 U7005 ( .B(n4788), .A(n3216), .Z(n4854) );
  CMX2X1 U7006 ( .A0(n4755), .A1(n4754), .S(n3213), .Z(n4878) );
  CMX2X1 U7007 ( .A0(n5150), .A1(n5217), .S(n3213), .Z(n5270) );
  CMX2X1 U7008 ( .A0(n5124), .A1(n5199), .S(n3207), .Z(n5261) );
  CMX2X1 U7009 ( .A0(n5116), .A1(n5195), .S(n3213), .Z(n5259) );
  CMX2X1 U7010 ( .A0(n5106), .A1(n5191), .S(n3199), .Z(n5257) );
  CMX2X1 U7011 ( .A0(n5101), .A1(n5188), .S(n3201), .Z(n5256) );
  CMX2X1 U7012 ( .A0(n4807), .A1(n4808), .S(n3209), .Z(n4873) );
  CAN2X1 U7013 ( .A(n5187), .B(n3203), .Z(n5255) );
  CAN2X1 U7014 ( .A(n4806), .B(n3216), .Z(n4908) );
  CAN2X1 U7015 ( .A(n4806), .B(n3203), .Z(n4872) );
  CAN2X1 U7016 ( .A(n5751), .B(n3213), .Z(n5817) );
  CAN2X1 U7017 ( .A(n6226), .B(n3210), .Z(n6327) );
  CAN2X1 U7018 ( .A(n6226), .B(n3199), .Z(n6292) );
  CAN2X1 U7019 ( .A(n5751), .B(n3214), .Z(n5853) );
  CMX2X1 U7020 ( .A0(n5131), .A1(n5203), .S(n3207), .Z(n5263) );
  CMX2X1 U7021 ( .A0(n13772), .A1(n13787), .S(n3790), .Z(n13800) );
  CND2X1 U7022 ( .A(n5134), .B(n3207), .Z(n5206) );
  CAN2X1 U7023 ( .A(n4804), .B(n3209), .Z(n4871) );
  CAN2X1 U7024 ( .A(n4775), .B(n3211), .Z(n4841) );
  CND2X1 U7025 ( .A(n5725), .B(n3205), .Z(n5791) );
  CND2X1 U7026 ( .A(n5720), .B(n3209), .Z(n5787) );
  CND2X1 U7027 ( .A(n5737), .B(n3211), .Z(n5803) );
  CND2X1 U7028 ( .A(n5746), .B(n3201), .Z(n5812) );
  CND2X1 U7029 ( .A(n5744), .B(n3215), .Z(n5810) );
  CND2X1 U7030 ( .A(n5735), .B(n3211), .Z(n5801) );
  CND2X1 U7031 ( .A(n5733), .B(n3199), .Z(n5799) );
  CND2X1 U7032 ( .A(n5731), .B(n3199), .Z(n5797) );
  CND2X1 U7033 ( .A(n5729), .B(n3207), .Z(n5795) );
  CND2X1 U7034 ( .A(n5718), .B(n3213), .Z(n5785) );
  CND2X1 U7035 ( .A(n6154), .B(n3207), .Z(n6228) );
  CND2X1 U7036 ( .A(n6158), .B(n3205), .Z(n6230) );
  CND2X1 U7037 ( .A(n5748), .B(n3215), .Z(n5814) );
  CND2X1 U7038 ( .A(n5155), .B(n3199), .Z(n5222) );
  CND2X1 U7039 ( .A(n6161), .B(n3215), .Z(n6232) );
  CND2X1 U7040 ( .A(n6167), .B(n3215), .Z(n6236) );
  CND2X1 U7041 ( .A(n6164), .B(n3215), .Z(n6234) );
  CND2X1 U7042 ( .A(n5140), .B(n3199), .Z(n5210) );
  CND2X1 U7043 ( .A(n5131), .B(n3207), .Z(n5204) );
  CND2X1 U7044 ( .A(n5727), .B(n3209), .Z(n5793) );
  CND2X1 U7045 ( .A(n5716), .B(n3201), .Z(n5782) );
  CND2X1 U7046 ( .A(n5695), .B(n3205), .Z(n5768) );
  CND2X1 U7047 ( .A(n5146), .B(n3205), .Z(n5216) );
  CND2X1 U7048 ( .A(n5143), .B(n3199), .Z(n5214) );
  CND2X1 U7049 ( .A(n5128), .B(n3213), .Z(n5202) );
  CND2X1 U7050 ( .A(n5116), .B(n3199), .Z(n5196) );
  CND2X1 U7051 ( .A(n5101), .B(n3201), .Z(n5189) );
  CND2X1 U7052 ( .A(n6173), .B(n3199), .Z(n6240) );
  CND2X1 U7053 ( .A(n6170), .B(n3203), .Z(n6238) );
  CND2X1 U7054 ( .A(n5710), .B(n3209), .Z(n5778) );
  CND2X1 U7055 ( .A(n5704), .B(n3215), .Z(n5774) );
  CND2X1 U7056 ( .A(n5248), .B(n3210), .Z(n5350) );
  CND2X1 U7057 ( .A(n5723), .B(n3199), .Z(n5789) );
  CND2X1 U7058 ( .A(n5713), .B(n3201), .Z(n5780) );
  CND2X1 U7059 ( .A(n5701), .B(n3207), .Z(n5772) );
  CND2X1 U7060 ( .A(n5698), .B(n3201), .Z(n5770) );
  CND2X1 U7061 ( .A(n5691), .B(n3207), .Z(n5766) );
  CND2X1 U7062 ( .A(n5687), .B(n3207), .Z(n5764) );
  CND2X1 U7063 ( .A(n5683), .B(n3215), .Z(n5761) );
  CND2X1 U7064 ( .A(n5675), .B(n3213), .Z(n5757) );
  CND2X1 U7065 ( .A(n5670), .B(n3199), .Z(n5755) );
  CND2X1 U7066 ( .A(n5665), .B(n3211), .Z(n5753) );
  CND2X1 U7067 ( .A(n5252), .B(n3212), .Z(n5354) );
  CND2X1 U7068 ( .A(n5137), .B(n3205), .Z(n5208) );
  CND2X1 U7069 ( .A(n5111), .B(n3209), .Z(n5194) );
  CND2X1 U7070 ( .A(n5106), .B(n3215), .Z(n5192) );
  CND2X1 U7071 ( .A(n4811), .B(n3207), .Z(n6512) );
  CND2X1 U7072 ( .A(n4809), .B(n3205), .Z(n6499) );
  CND2X1 U7073 ( .A(n4807), .B(n3203), .Z(n6486) );
  CND2X1 U7074 ( .A(n5679), .B(n3205), .Z(n5759) );
  CND2X1 U7075 ( .A(n5773), .B(n3216), .Z(n5875) );
  CND2X1 U7076 ( .A(n5777), .B(n3204), .Z(n5880) );
  CND2X1 U7077 ( .A(n5769), .B(n3212), .Z(n5871) );
  CND2X1 U7078 ( .A(n5765), .B(n3204), .Z(n5867) );
  CND2X1 U7079 ( .A(n5760), .B(n3200), .Z(n5863) );
  CND2X1 U7080 ( .A(n5752), .B(n3206), .Z(n5854) );
  CND2X1 U7081 ( .A(n4812), .B(n3216), .Z(n4914) );
  CND2X1 U7082 ( .A(n5779), .B(n3208), .Z(n5882) );
  CND2X1 U7083 ( .A(n5756), .B(n3206), .Z(n5859) );
  CND2X1 U7084 ( .A(n5754), .B(n3210), .Z(n5857) );
  CND2X1 U7085 ( .A(n5758), .B(n3212), .Z(n5861) );
  CND2X1 U7086 ( .A(n6239), .B(n3206), .Z(n6341) );
  CND2X1 U7087 ( .A(n6237), .B(n3202), .Z(n6339) );
  CND2X1 U7088 ( .A(n6227), .B(n3214), .Z(n6328) );
  CND2X1 U7089 ( .A(n5767), .B(n3212), .Z(n5869) );
  CND2X1 U7090 ( .A(n5225), .B(n3210), .Z(n5327) );
  CND2X1 U7091 ( .A(n6229), .B(n3202), .Z(n6330) );
  CND2X1 U7092 ( .A(n5238), .B(n3202), .Z(n5339) );
  CND2X1 U7093 ( .A(n5781), .B(n3208), .Z(n5884) );
  CND2X1 U7094 ( .A(n5236), .B(n3206), .Z(n5337) );
  CND2X1 U7095 ( .A(n6231), .B(n3214), .Z(n6332) );
  CND2X1 U7096 ( .A(n5813), .B(n3200), .Z(n5915) );
  CND2X1 U7097 ( .A(n5234), .B(n3212), .Z(n5335) );
  CND2X1 U7098 ( .A(n5231), .B(n3208), .Z(n5333) );
  CND2X1 U7099 ( .A(n5229), .B(n3204), .Z(n5331) );
  CND2X1 U7100 ( .A(n5227), .B(n3216), .Z(n5329) );
  CND2X1 U7101 ( .A(n5221), .B(n3200), .Z(n5322) );
  CND2X1 U7102 ( .A(n6233), .B(n3216), .Z(n6334) );
  CND2X1 U7103 ( .A(n6235), .B(n3210), .Z(n6336) );
  CND2X1 U7104 ( .A(n5815), .B(n3216), .Z(n5917) );
  CND2X1 U7105 ( .A(n5811), .B(n3206), .Z(n5913) );
  CND2X1 U7106 ( .A(n5809), .B(n3208), .Z(n5911) );
  CND2X1 U7107 ( .A(n5807), .B(n3200), .Z(n5909) );
  CND2X1 U7108 ( .A(n5805), .B(n3204), .Z(n5907) );
  CND2X1 U7109 ( .A(n5802), .B(n3202), .Z(n5905) );
  CND2X1 U7110 ( .A(n5800), .B(n3210), .Z(n5903) );
  CND2X1 U7111 ( .A(n5798), .B(n3216), .Z(n5901) );
  CND2X1 U7112 ( .A(n5796), .B(n3206), .Z(n5899) );
  CND2X1 U7113 ( .A(n5794), .B(n3210), .Z(n5896) );
  CND2X1 U7114 ( .A(n5790), .B(n3216), .Z(n5892) );
  CND2X1 U7115 ( .A(n5786), .B(n3202), .Z(n5888) );
  CND2X1 U7116 ( .A(n5784), .B(n3214), .Z(n5886) );
  CND2X1 U7117 ( .A(n5775), .B(n3208), .Z(n5878) );
  CND2X1 U7118 ( .A(n5771), .B(n3204), .Z(n5873) );
  CND2X1 U7119 ( .A(n5763), .B(n3200), .Z(n5865) );
  CND2X1 U7120 ( .A(n5244), .B(n3204), .Z(n5345) );
  CND2X1 U7121 ( .A(n5250), .B(n3214), .Z(n5352) );
  CND2X1 U7122 ( .A(n5246), .B(n3216), .Z(n5348) );
  CND2X1 U7123 ( .A(n5242), .B(n3206), .Z(n5343) );
  CND2X1 U7124 ( .A(n5240), .B(n3202), .Z(n5341) );
  CIVX2 U7125 ( .A(n4193), .Z(n3750) );
  CNR2X1 U7126 ( .A(n3511), .B(n6575), .Z(N3098) );
  CNR2X1 U7127 ( .A(n3510), .B(n6576), .Z(N3099) );
  COR2X1 U7128 ( .A(n3692), .B(n3682), .Z(n2105) );
  CMXI2X1 U7129 ( .A0(n13741), .A1(n15076), .S(n3804), .Z(n13743) );
  CMXI2X1 U7130 ( .A0(n13404), .A1(n14742), .S(n3804), .Z(n13406) );
  CMX2X1 U7131 ( .A0(n3745), .A1(n4801), .S(n3211), .Z(n4906) );
  CMXI2X1 U7132 ( .A0(n10669), .A1(n12005), .S(n3803), .Z(n10671) );
  CEOX1 U7133 ( .A(N3109), .B(n3266), .Z(N6231) );
  CNR2X1 U7134 ( .A(N3108), .B(\r349/carry [8]), .Z(n3266) );
  CNR2IX1 U7135 ( .B(n4802), .A(n3208), .Z(n4869) );
  CNR2IX1 U7136 ( .B(n4798), .A(n3214), .Z(n4864) );
  CNR2IX1 U7137 ( .B(n4770), .A(n3215), .Z(n4836) );
  CNR2IX1 U7138 ( .B(n6214), .A(n3209), .Z(n6281) );
  CNR2IX1 U7139 ( .B(n6212), .A(n3215), .Z(n6279) );
  CNR2IX1 U7140 ( .B(n6210), .A(n3203), .Z(n6277) );
  CNR2X1 U7141 ( .A(n3826), .B(n5389), .Z(N431) );
  CNR2X1 U7142 ( .A(n3764), .B(n5053), .Z(n5137) );
  CNR2X1 U7143 ( .A(n3765), .B(n5045), .Z(n5134) );
  CNR2X1 U7144 ( .A(n5038), .B(n3765), .Z(n5131) );
  CNR2X1 U7145 ( .A(n5003), .B(n3765), .Z(n5111) );
  CNR2X1 U7146 ( .A(n4989), .B(n3765), .Z(n5101) );
  CNR2X1 U7147 ( .A(n4739), .B(n3764), .Z(n4807) );
  CNR2X1 U7148 ( .A(n3763), .B(n5060), .Z(n5140) );
  CNR2X1 U7149 ( .A(n3762), .B(n5095), .Z(n5155) );
  CNR2X1 U7150 ( .A(n6123), .B(n3766), .Z(n6173) );
  CNR2X1 U7151 ( .A(n6119), .B(n3763), .Z(n6170) );
  CNR2X1 U7152 ( .A(n6115), .B(n3766), .Z(n6167) );
  CNR2X1 U7153 ( .A(n6111), .B(n3763), .Z(n6164) );
  CNR2X1 U7154 ( .A(n6107), .B(n3762), .Z(n6161) );
  CNR2X1 U7155 ( .A(n6103), .B(n3762), .Z(n6158) );
  CNR2X1 U7156 ( .A(n6099), .B(n3762), .Z(n6154) );
  CNR2X1 U7157 ( .A(n3763), .B(n5637), .Z(n5710) );
  CNR2X1 U7158 ( .A(n3766), .B(n5630), .Z(n5707) );
  CNR2X1 U7159 ( .A(n3766), .B(n5623), .Z(n5704) );
  CNR2X1 U7160 ( .A(n3766), .B(n5659), .Z(n5718) );
  CNR2X1 U7161 ( .A(n3764), .B(n5652), .Z(n5716) );
  CNR2X1 U7162 ( .A(n3762), .B(n5645), .Z(n5713) );
  CNR2X1 U7163 ( .A(n3765), .B(n5616), .Z(n5701) );
  CNR2X1 U7164 ( .A(n3764), .B(n5609), .Z(n5698) );
  CNR2X1 U7165 ( .A(n5602), .B(n3762), .Z(n5695) );
  CNR2X1 U7166 ( .A(n5595), .B(n3763), .Z(n5691) );
  CNR2X1 U7167 ( .A(n5588), .B(n3764), .Z(n5687) );
  CNR2X1 U7168 ( .A(n5581), .B(n3766), .Z(n5683) );
  CNR2X1 U7169 ( .A(n5565), .B(n3766), .Z(n5675) );
  CNR2X1 U7170 ( .A(n5558), .B(n3763), .Z(n5670) );
  CNR2X1 U7171 ( .A(n5551), .B(n3766), .Z(n5665) );
  CNR2X1 U7172 ( .A(n4744), .B(n3764), .Z(n4809) );
  CNR2X1 U7173 ( .A(n5574), .B(n3765), .Z(n5679) );
  CNR2X1 U7174 ( .A(n5168), .B(n3761), .Z(n5236) );
  CNR2X1 U7175 ( .A(n5164), .B(n3761), .Z(n5231) );
  CNR2X1 U7176 ( .A(n5158), .B(n3760), .Z(n5225) );
  CNR2X1 U7177 ( .A(n5166), .B(n3760), .Z(n5234) );
  CNR2X1 U7178 ( .A(n5154), .B(n3760), .Z(n5221) );
  CNR2X1 U7179 ( .A(n5749), .B(n3759), .Z(n5815) );
  CNR2X1 U7180 ( .A(n5743), .B(n3761), .Z(n5809) );
  CNR2X1 U7181 ( .A(n5740), .B(n3761), .Z(n5807) );
  CNR2X1 U7182 ( .A(n5738), .B(n3758), .Z(n5805) );
  CNR2X1 U7183 ( .A(n5736), .B(n3760), .Z(n5802) );
  CNR2X1 U7184 ( .A(n5734), .B(n3759), .Z(n5800) );
  CNR2X1 U7185 ( .A(n5732), .B(n3758), .Z(n5798) );
  CNR2X1 U7186 ( .A(n5730), .B(n3760), .Z(n5796) );
  CNR2X1 U7187 ( .A(n5728), .B(n3758), .Z(n5794) );
  CNR2X1 U7188 ( .A(n5724), .B(n3761), .Z(n5790) );
  CNR2X1 U7189 ( .A(n5719), .B(n3761), .Z(n5786) );
  CNR2X1 U7190 ( .A(n5717), .B(n3758), .Z(n5784) );
  CNR2X1 U7191 ( .A(n5185), .B(n3759), .Z(n5252) );
  CNR2X1 U7192 ( .A(n5183), .B(n3759), .Z(n5250) );
  CNR2X1 U7193 ( .A(n5179), .B(n3759), .Z(n5246) );
  CNR2X1 U7194 ( .A(n5177), .B(n3758), .Z(n5244) );
  CNR2X1 U7195 ( .A(n5173), .B(n3760), .Z(n5240) );
  CND2X1 U7196 ( .A(n3727), .B(n5280), .Z(n5382) );
  CNR2X1 U7197 ( .A(n4697), .B(n3764), .Z(n4755) );
  CNR2X1 U7198 ( .A(n3763), .B(n4669), .Z(n4773) );
  CNR2X1 U7199 ( .A(n4707), .B(n3762), .Z(n4759) );
  CNR2X1 U7200 ( .A(n3766), .B(n6144), .Z(n6188) );
  CNR2X1 U7201 ( .A(n4693), .B(n3765), .Z(n4753) );
  CNR2X1 U7202 ( .A(n3766), .B(n4735), .Z(n4771) );
  CNR2X1 U7203 ( .A(n3765), .B(n6150), .Z(n6192) );
  CNR2X1 U7204 ( .A(n3762), .B(n6141), .Z(n6186) );
  CNR2X1 U7205 ( .A(n3762), .B(n6138), .Z(n6184) );
  CNR2X1 U7206 ( .A(n3762), .B(n6135), .Z(n6181) );
  CNR2X1 U7207 ( .A(n3764), .B(n6132), .Z(n6179) );
  CNR2X1 U7208 ( .A(n3765), .B(n6129), .Z(n6177) );
  CNR2X1 U7209 ( .A(n6126), .B(n3764), .Z(n6175) );
  CNR2X1 U7210 ( .A(n6163), .B(n3759), .Z(n6199) );
  CNR2X1 U7211 ( .A(n6166), .B(n3758), .Z(n6201) );
  CNR2X1 U7212 ( .A(n6151), .B(n3759), .Z(n6191) );
  CNR2X1 U7213 ( .A(n6160), .B(n3758), .Z(n6197) );
  CNR2X1 U7214 ( .A(n6157), .B(n3760), .Z(n6195) );
  CNR2X1 U7215 ( .A(n4568), .B(n3760), .Z(n6216) );
  CNR2X1 U7216 ( .A(n4532), .B(n3760), .Z(n6210) );
  CNR2X1 U7217 ( .A(n4531), .B(n3761), .Z(n6208) );
  CNR2X1 U7218 ( .A(n4692), .B(n3760), .Z(n4782) );
  CNR2X1 U7219 ( .A(n4668), .B(n3759), .Z(n4772) );
  CNR2X1 U7220 ( .A(n4571), .B(n3761), .Z(n6222) );
  CNR2X1 U7221 ( .A(n4910), .B(n4207), .Z(n4913) );
  CNR2X1 U7222 ( .A(n6030), .B(n4208), .Z(n6034) );
  CNR2X1 U7223 ( .A(n5467), .B(n4207), .Z(n5471) );
  CNR2X1 U7224 ( .A(n4566), .B(n4210), .Z(n4604) );
  CND2X1 U7225 ( .A(n3725), .B(n5841), .Z(n5944) );
  CND2X1 U7226 ( .A(n6293), .B(n3740), .Z(n6466) );
  CND2X1 U7227 ( .A(n3730), .B(n6293), .Z(n6394) );
  CND2X1 U7228 ( .A(n3723), .B(n6299), .Z(n6402) );
  CND2X1 U7229 ( .A(n5841), .B(n3735), .Z(n6015) );
  CND2X1 U7230 ( .A(n5840), .B(n3734), .Z(n6014) );
  CND2X1 U7231 ( .A(n3725), .B(n5840), .Z(n5943) );
  CND2X1 U7232 ( .A(n6326), .B(n3737), .Z(n6503) );
  CND2X1 U7233 ( .A(n6299), .B(n3736), .Z(n6472) );
  CND2X1 U7234 ( .A(n3725), .B(n5842), .Z(n5945) );
  CND2X1 U7235 ( .A(n3724), .B(n6301), .Z(n6403) );
  CND2X1 U7236 ( .A(n3722), .B(n6298), .Z(n6401) );
  CND2X1 U7237 ( .A(n6298), .B(n3735), .Z(n6471) );
  CND2X1 U7238 ( .A(n5848), .B(n3733), .Z(n6021) );
  CND2X1 U7239 ( .A(n5831), .B(n3735), .Z(n6005) );
  CND2X1 U7240 ( .A(n5828), .B(n3737), .Z(n6002) );
  CND2X1 U7241 ( .A(n3726), .B(n5846), .Z(n5947) );
  CND2X1 U7242 ( .A(n3728), .B(n5831), .Z(n5934) );
  CND2X1 U7243 ( .A(n3727), .B(n5828), .Z(n5931) );
  CND2X1 U7244 ( .A(n6309), .B(n3738), .Z(n6482) );
  CND2X1 U7245 ( .A(n6303), .B(n3733), .Z(n6476) );
  CND2X1 U7246 ( .A(n6301), .B(n3734), .Z(n6473) );
  CND2X1 U7247 ( .A(n5851), .B(n3731), .Z(n6024) );
  CND2X1 U7248 ( .A(n6310), .B(n3740), .Z(n6483) );
  CND2X1 U7249 ( .A(n6307), .B(n3731), .Z(n6480) );
  CND2X1 U7250 ( .A(n6306), .B(n3733), .Z(n6479) );
  CND2X1 U7251 ( .A(n6304), .B(n3735), .Z(n6477) );
  CND2X1 U7252 ( .A(n3726), .B(n6326), .Z(n6428) );
  CND2X1 U7253 ( .A(n3726), .B(n6310), .Z(n6413) );
  CND2X1 U7254 ( .A(n3722), .B(n6309), .Z(n6412) );
  CND2X1 U7255 ( .A(n3727), .B(n6304), .Z(n6406) );
  CND2X1 U7256 ( .A(n3727), .B(n6303), .Z(n6405) );
  CND2X1 U7257 ( .A(n5852), .B(n3738), .Z(n6025) );
  CND2X1 U7258 ( .A(n5846), .B(n3734), .Z(n6018) );
  CND2X1 U7259 ( .A(n5842), .B(n3732), .Z(n6016) );
  CND2X1 U7260 ( .A(n5839), .B(n3732), .Z(n6013) );
  CND2X1 U7261 ( .A(n5836), .B(n3740), .Z(n6010) );
  CND2X1 U7262 ( .A(n5834), .B(n3736), .Z(n6007) );
  CND2X1 U7263 ( .A(n3722), .B(n5852), .Z(n5954) );
  CND2X1 U7264 ( .A(n3729), .B(n5836), .Z(n5938) );
  CND2X1 U7265 ( .A(n3726), .B(n5834), .Z(n5936) );
  CND2X1 U7266 ( .A(n3723), .B(n5820), .Z(n5923) );
  CND2X1 U7267 ( .A(n6294), .B(n3733), .Z(n6467) );
  CND2X1 U7268 ( .A(n6325), .B(n3733), .Z(n6502) );
  CND2X1 U7269 ( .A(n6318), .B(n3740), .Z(n6493) );
  CND2X1 U7270 ( .A(n3726), .B(n6307), .Z(n6410) );
  CND2X1 U7271 ( .A(n3724), .B(n6306), .Z(n6408) );
  CND2X1 U7272 ( .A(n3723), .B(n6294), .Z(n6395) );
  CND2X1 U7273 ( .A(n5833), .B(n3739), .Z(n6006) );
  CND2X1 U7274 ( .A(n5827), .B(n3740), .Z(n6001) );
  CND2X1 U7275 ( .A(n5818), .B(n3731), .Z(n5992) );
  CND2X1 U7276 ( .A(n3726), .B(n5850), .Z(n5951) );
  CND2X1 U7277 ( .A(n3726), .B(n5849), .Z(n5950) );
  CND2X1 U7278 ( .A(n3728), .B(n5845), .Z(n5946) );
  CND2X1 U7279 ( .A(n3729), .B(n5833), .Z(n5935) );
  CND2X1 U7280 ( .A(n3730), .B(n5827), .Z(n5929) );
  CND2X1 U7281 ( .A(n3730), .B(n5818), .Z(n5921) );
  CND2X1 U7282 ( .A(n5255), .B(n3740), .Z(n5427) );
  CND2X1 U7283 ( .A(n3723), .B(n4887), .Z(n4767) );
  CND2X1 U7284 ( .A(n3726), .B(n4886), .Z(n4766) );
  CND2X1 U7285 ( .A(n3725), .B(n4885), .Z(n4763) );
  CND2X1 U7286 ( .A(n3724), .B(n4884), .Z(n4762) );
  CND2X1 U7287 ( .A(n3725), .B(n4882), .Z(n6398) );
  CND2X1 U7288 ( .A(n3727), .B(n4878), .Z(n5986) );
  CND2X1 U7289 ( .A(n3730), .B(n4877), .Z(n5844) );
  CND2X1 U7290 ( .A(n3727), .B(n4875), .Z(n5374) );
  CND2X1 U7291 ( .A(n3730), .B(n4874), .Z(n5212) );
  CND2X1 U7292 ( .A(n6324), .B(n3734), .Z(n6498) );
  CND2X1 U7293 ( .A(n6308), .B(n3739), .Z(n6481) );
  CND2X1 U7294 ( .A(n6302), .B(n3737), .Z(n6474) );
  CND2X1 U7295 ( .A(n6323), .B(n3737), .Z(n6497) );
  CND2X1 U7296 ( .A(n3728), .B(n5286), .Z(n5389) );
  CND2X1 U7297 ( .A(n6321), .B(n3731), .Z(n6496) );
  CND2X1 U7298 ( .A(n6320), .B(n3733), .Z(n6495) );
  CND2X1 U7299 ( .A(n6319), .B(n3738), .Z(n6494) );
  CND2X1 U7300 ( .A(n6316), .B(n3734), .Z(n6491) );
  CND2X1 U7301 ( .A(n6315), .B(n3733), .Z(n6490) );
  CND2X1 U7302 ( .A(n6314), .B(n3736), .Z(n6489) );
  CND2X1 U7303 ( .A(n6313), .B(n3736), .Z(n6485) );
  CND2X1 U7304 ( .A(n6312), .B(n3740), .Z(n6484) );
  CND2X1 U7305 ( .A(n6305), .B(n3737), .Z(n6478) );
  CND2X1 U7306 ( .A(n6297), .B(n3731), .Z(n6470) );
  CND2X1 U7307 ( .A(n6296), .B(n3737), .Z(n6469) );
  CND2X1 U7308 ( .A(n6295), .B(n3735), .Z(n6468) );
  CND2X1 U7309 ( .A(n3724), .B(n6325), .Z(n6427) );
  CND2X1 U7310 ( .A(n3724), .B(n6324), .Z(n6426) );
  CND2X1 U7311 ( .A(n3726), .B(n6323), .Z(n6425) );
  CND2X1 U7312 ( .A(n3727), .B(n6321), .Z(n6424) );
  CND2X1 U7313 ( .A(n3724), .B(n6320), .Z(n6423) );
  CND2X1 U7314 ( .A(n3722), .B(n6319), .Z(n6422) );
  CND2X1 U7315 ( .A(n3723), .B(n6318), .Z(n6421) );
  CND2X1 U7316 ( .A(n3730), .B(n6317), .Z(n6419) );
  CND2X1 U7317 ( .A(n3729), .B(n6316), .Z(n6418) );
  CND2X1 U7318 ( .A(n3724), .B(n6315), .Z(n6417) );
  CND2X1 U7319 ( .A(n3729), .B(n6314), .Z(n6416) );
  CND2X1 U7320 ( .A(n3725), .B(n6313), .Z(n6415) );
  CND2X1 U7321 ( .A(n3728), .B(n6312), .Z(n6414) );
  CND2X1 U7322 ( .A(n3723), .B(n6308), .Z(n6411) );
  CND2X1 U7323 ( .A(n3722), .B(n6305), .Z(n6407) );
  CND2X1 U7324 ( .A(n3724), .B(n6302), .Z(n6404) );
  CND2X1 U7325 ( .A(n3723), .B(n6297), .Z(n6400) );
  CND2X1 U7326 ( .A(n3728), .B(n6296), .Z(n6399) );
  CND2X1 U7327 ( .A(n3730), .B(n6295), .Z(n6396) );
  CND2X1 U7328 ( .A(n5845), .B(n3740), .Z(n6017) );
  CND2X1 U7329 ( .A(n5838), .B(n3737), .Z(n6012) );
  CND2X1 U7330 ( .A(n5837), .B(n3734), .Z(n6011) );
  CND2X1 U7331 ( .A(n5826), .B(n3740), .Z(n6000) );
  CND2X1 U7332 ( .A(n5825), .B(n3732), .Z(n5999) );
  CND2X1 U7333 ( .A(n5824), .B(n3738), .Z(n5998) );
  CND2X1 U7334 ( .A(n5822), .B(n3739), .Z(n5995) );
  CND2X1 U7335 ( .A(n5820), .B(n3731), .Z(n5994) );
  CND2X1 U7336 ( .A(n5819), .B(n3732), .Z(n5993) );
  CND2X1 U7337 ( .A(n3724), .B(n5851), .Z(n5953) );
  CND2X1 U7338 ( .A(n3722), .B(n5848), .Z(n5949) );
  CND2X1 U7339 ( .A(n3727), .B(n5839), .Z(n5942) );
  CND2X1 U7340 ( .A(n3726), .B(n5838), .Z(n5940) );
  CND2X1 U7341 ( .A(n3722), .B(n5837), .Z(n5939) );
  CND2X1 U7342 ( .A(n3730), .B(n5826), .Z(n5928) );
  CND2X1 U7343 ( .A(n3726), .B(n5825), .Z(n5927) );
  CND2X1 U7344 ( .A(n3728), .B(n5824), .Z(n5926) );
  CND2X1 U7345 ( .A(n3725), .B(n5819), .Z(n5922) );
  CND2X1 U7346 ( .A(n5289), .B(n3732), .Z(n5461) );
  CND2X1 U7347 ( .A(n5284), .B(n3732), .Z(n5457) );
  CND2X1 U7348 ( .A(n5288), .B(n3736), .Z(n5460) );
  CND2X1 U7349 ( .A(n5283), .B(n3735), .Z(n5456) );
  CND2X1 U7350 ( .A(n5282), .B(n3734), .Z(n5455) );
  CND2X1 U7351 ( .A(n5281), .B(n3731), .Z(n5454) );
  CND2X1 U7352 ( .A(n5280), .B(n3733), .Z(n5453) );
  CND2X1 U7353 ( .A(n5279), .B(n3732), .Z(n5452) );
  CND2X1 U7354 ( .A(n5278), .B(n3733), .Z(n5450) );
  CND2X1 U7355 ( .A(n5277), .B(n3734), .Z(n5449) );
  CND2X1 U7356 ( .A(n5274), .B(n3737), .Z(n5447) );
  CND2X1 U7357 ( .A(n5272), .B(n3735), .Z(n5445) );
  CND2X1 U7358 ( .A(n5271), .B(n3734), .Z(n5444) );
  CND2X1 U7359 ( .A(n5270), .B(n3735), .Z(n5443) );
  CND2X1 U7360 ( .A(n5269), .B(n3731), .Z(n5442) );
  CND2X1 U7361 ( .A(n5268), .B(n3737), .Z(n5441) );
  CND2X1 U7362 ( .A(n5266), .B(n3736), .Z(n5438) );
  CND2X1 U7363 ( .A(n5264), .B(n3736), .Z(n5437) );
  CND2X1 U7364 ( .A(n5262), .B(n3739), .Z(n5435) );
  CND2X1 U7365 ( .A(n5261), .B(n3735), .Z(n5434) );
  CND2X1 U7366 ( .A(n5260), .B(n3738), .Z(n5433) );
  CND2X1 U7367 ( .A(n5259), .B(n3739), .Z(n5432) );
  CND2X1 U7368 ( .A(n5258), .B(n3732), .Z(n5431) );
  CND2X1 U7369 ( .A(n5257), .B(n3734), .Z(n5430) );
  CND2X1 U7370 ( .A(n5256), .B(n3738), .Z(n5428) );
  CND2X1 U7371 ( .A(n5290), .B(n3726), .Z(n5392) );
  CND2X1 U7372 ( .A(n3723), .B(n5289), .Z(n5391) );
  CND2X1 U7373 ( .A(n3730), .B(n5288), .Z(n5390) );
  CND2X1 U7374 ( .A(n3723), .B(n5284), .Z(n5387) );
  CND2X1 U7375 ( .A(n3725), .B(n5283), .Z(n5386) );
  CND2X1 U7376 ( .A(n3723), .B(n5282), .Z(n5384) );
  CND2X1 U7377 ( .A(n3724), .B(n5281), .Z(n5383) );
  CND2X1 U7378 ( .A(n3723), .B(n5279), .Z(n5381) );
  CND2X1 U7379 ( .A(n3729), .B(n5278), .Z(n5380) );
  CND2X1 U7380 ( .A(n3730), .B(n5277), .Z(n5379) );
  CND2X1 U7381 ( .A(n3726), .B(n5274), .Z(n5377) );
  CND2X1 U7382 ( .A(n3729), .B(n5272), .Z(n5375) );
  CND2X1 U7383 ( .A(n3728), .B(n5271), .Z(n5372) );
  CND2X1 U7384 ( .A(n3727), .B(n5270), .Z(n5371) );
  CND2X1 U7385 ( .A(n3725), .B(n5269), .Z(n5370) );
  CND2X1 U7386 ( .A(n3729), .B(n5268), .Z(n5369) );
  CND2X1 U7387 ( .A(n3726), .B(n5267), .Z(n5368) );
  CND2X1 U7388 ( .A(n3729), .B(n5266), .Z(n5367) );
  CND2X1 U7389 ( .A(n3721), .B(n5264), .Z(n5366) );
  CND2X1 U7390 ( .A(n3730), .B(n5262), .Z(n5364) );
  CND2X1 U7391 ( .A(n3721), .B(n5261), .Z(n5363) );
  CND2X1 U7392 ( .A(n3723), .B(n5259), .Z(n5360) );
  CND2X1 U7393 ( .A(n3726), .B(n5258), .Z(n5359) );
  CND2X1 U7394 ( .A(n3722), .B(n5257), .Z(n5358) );
  CND2X1 U7395 ( .A(n3728), .B(n5256), .Z(n5357) );
  CND2X1 U7396 ( .A(n4908), .B(n3737), .Z(n6475) );
  CND2X1 U7397 ( .A(n4907), .B(n3731), .Z(n6464) );
  CND2X1 U7398 ( .A(n4906), .B(n3736), .Z(n6453) );
  CND2X1 U7399 ( .A(n4905), .B(n3731), .Z(n6442) );
  CND2X1 U7400 ( .A(n4904), .B(n3733), .Z(n6431) );
  CND2X1 U7401 ( .A(n4902), .B(n3733), .Z(n6420) );
  CND2X1 U7402 ( .A(n4901), .B(n3731), .Z(n6409) );
  CND2X1 U7403 ( .A(n4899), .B(n3740), .Z(n6380) );
  CND2X1 U7404 ( .A(n4898), .B(n3732), .Z(n6359) );
  CND2X1 U7405 ( .A(n4897), .B(n3732), .Z(n6338) );
  CND2X1 U7406 ( .A(n4896), .B(n3739), .Z(n6322) );
  CND2X1 U7407 ( .A(n4895), .B(n3736), .Z(n6311) );
  CND2X1 U7408 ( .A(n4894), .B(n3738), .Z(n6300) );
  CND2X1 U7409 ( .A(n4893), .B(n3734), .Z(n6287) );
  CND2X1 U7410 ( .A(n4891), .B(n3732), .Z(n6266) );
  CND2X1 U7411 ( .A(n4890), .B(n3736), .Z(n6245) );
  CND2X1 U7412 ( .A(n4889), .B(n3737), .Z(n6224) );
  CND2X1 U7413 ( .A(n4878), .B(n3739), .Z(n5997) );
  CND2X1 U7414 ( .A(n4877), .B(n3740), .Z(n5985) );
  CND2X1 U7415 ( .A(n4876), .B(n3739), .Z(n5974) );
  CND2X1 U7416 ( .A(n4875), .B(n3732), .Z(n5963) );
  CND2X1 U7417 ( .A(n4874), .B(n3735), .Z(n5952) );
  CND2X1 U7418 ( .A(n4873), .B(n3739), .Z(n5941) );
  CND2X1 U7419 ( .A(n4872), .B(n3732), .Z(n5930) );
  CND2X1 U7420 ( .A(n4908), .B(n3730), .Z(n5265) );
  CND2X1 U7421 ( .A(n3729), .B(n4907), .Z(n5254) );
  CND2X1 U7422 ( .A(n3723), .B(n4906), .Z(n5233) );
  CND2X1 U7423 ( .A(n3728), .B(n4905), .Z(n5211) );
  CND2X1 U7424 ( .A(n3730), .B(n4904), .Z(n5190) );
  CND2X1 U7425 ( .A(n3730), .B(n4902), .Z(n5170) );
  CND2X1 U7426 ( .A(n3725), .B(n4901), .Z(n5147) );
  CND2X1 U7427 ( .A(n3729), .B(n4899), .Z(n5047) );
  CND2X1 U7428 ( .A(n3727), .B(n4898), .Z(n4977) );
  CND2X1 U7429 ( .A(n3724), .B(n4897), .Z(n4922) );
  CND2X1 U7430 ( .A(n3728), .B(n4896), .Z(n4903) );
  CND2X1 U7431 ( .A(n3729), .B(n4895), .Z(n4892) );
  CND2X1 U7432 ( .A(n3722), .B(n4894), .Z(n4880) );
  CND2X1 U7433 ( .A(n3729), .B(n4893), .Z(n4867) );
  CND2X1 U7434 ( .A(n3727), .B(n4891), .Z(n4846) );
  CND2X1 U7435 ( .A(n3725), .B(n4890), .Z(n4825) );
  CND2X1 U7436 ( .A(n3725), .B(n4889), .Z(n4805) );
  CND2X1 U7437 ( .A(n3730), .B(n4873), .Z(n4881) );
  CND2X1 U7438 ( .A(n4872), .B(n3725), .Z(n4738) );
  CND2X1 U7439 ( .A(n6327), .B(n3736), .Z(n6504) );
  CND2X1 U7440 ( .A(n6292), .B(n3740), .Z(n6465) );
  CND2X1 U7441 ( .A(n6327), .B(n3727), .Z(n6429) );
  CND2X1 U7442 ( .A(n6292), .B(n3727), .Z(n6393) );
  CND2X1 U7443 ( .A(n5853), .B(n3739), .Z(n6026) );
  CND2X1 U7444 ( .A(n5847), .B(n3739), .Z(n6020) );
  CND2X1 U7445 ( .A(n5835), .B(n3738), .Z(n6009) );
  CND2X1 U7446 ( .A(n5830), .B(n3737), .Z(n6004) );
  CND2X1 U7447 ( .A(n5829), .B(n3738), .Z(n6003) );
  CND2X1 U7448 ( .A(n5853), .B(n3729), .Z(n5955) );
  CND2X1 U7449 ( .A(n3722), .B(n5847), .Z(n5948) );
  CND2X1 U7450 ( .A(n3729), .B(n5835), .Z(n5937) );
  CND2X1 U7451 ( .A(n3724), .B(n5830), .Z(n5933) );
  CND2X1 U7452 ( .A(n3730), .B(n5829), .Z(n5932) );
  CND2X1 U7453 ( .A(n3727), .B(n5822), .Z(n5924) );
  CNR2X1 U7454 ( .A(n5024), .B(n3764), .Z(n5124) );
  CND2X1 U7455 ( .A(n3730), .B(n4883), .Z(n6515) );
  CNR2X1 U7456 ( .A(n5017), .B(n3765), .Z(n5120) );
  CND2X1 U7457 ( .A(n5286), .B(n3736), .Z(n5459) );
  CND2X1 U7458 ( .A(n5273), .B(n3740), .Z(n5446) );
  CND2X1 U7459 ( .A(n5267), .B(n3733), .Z(n5439) );
  CND2X1 U7460 ( .A(n3723), .B(n5273), .Z(n5376) );
  CND2X1 U7461 ( .A(n3727), .B(n5260), .Z(n5361) );
  CIVX2 U7462 ( .A(n4298), .Z(n4267) );
  CIVX2 U7463 ( .A(n4299), .Z(n4270) );
  CIVX2 U7464 ( .A(n4299), .Z(n4272) );
  CMX2X1 U7465 ( .A0(n5111), .A1(n5193), .S(n3211), .Z(n5258) );
  CND2X1 U7466 ( .A(n4969), .B(n3894), .Z(n5024) );
  CND2X1 U7467 ( .A(n4945), .B(n3893), .Z(n4996) );
  CND2X1 U7468 ( .A(n5144), .B(n4222), .Z(n5181) );
  CNIVX1 U7469 ( .A(n4437), .Z(n4217) );
  CNIVX1 U7470 ( .A(n4437), .Z(n4218) );
  CNIVX1 U7471 ( .A(n4437), .Z(n4219) );
  CNIVX1 U7472 ( .A(n4437), .Z(n4215) );
  CND2X1 U7473 ( .A(n5849), .B(n3733), .Z(n6022) );
  CND2X1 U7474 ( .A(n6317), .B(n3737), .Z(n6492) );
  CND2X1 U7475 ( .A(n5850), .B(n3734), .Z(n6023) );
  CND2X1 U7476 ( .A(n5817), .B(n3735), .Z(n5991) );
  CND2X1 U7477 ( .A(n5817), .B(n3730), .Z(n5920) );
  CND2X1 U7478 ( .A(n6258), .B(n3736), .Z(n6361) );
  CND2X1 U7479 ( .A(n6260), .B(n3732), .Z(n6363) );
  CND2X1 U7480 ( .A(n6243), .B(n3732), .Z(n6346) );
  CND2X1 U7481 ( .A(n6241), .B(n3734), .Z(n6344) );
  CND2X1 U7482 ( .A(n6264), .B(n3738), .Z(n6367) );
  CND2X1 U7483 ( .A(n6256), .B(n3734), .Z(n6358) );
  CND2X1 U7484 ( .A(n6267), .B(n3735), .Z(n6369) );
  CND2X1 U7485 ( .A(n6262), .B(n3736), .Z(n6365) );
  CND2X1 U7486 ( .A(n6254), .B(n3737), .Z(n6356) );
  CND2X1 U7487 ( .A(n6271), .B(n3733), .Z(n6373) );
  CND2X1 U7488 ( .A(n6269), .B(n3731), .Z(n6371) );
  CND2X1 U7489 ( .A(n6285), .B(n3731), .Z(n6388) );
  CND2X1 U7490 ( .A(n6283), .B(n3735), .Z(n6386) );
  CND2X1 U7491 ( .A(n6281), .B(n3733), .Z(n6384) );
  CND2X1 U7492 ( .A(n6279), .B(n3740), .Z(n6382) );
  CND2X1 U7493 ( .A(n6277), .B(n3734), .Z(n6379) );
  CND2X1 U7494 ( .A(n6275), .B(n3739), .Z(n6377) );
  CND2X1 U7495 ( .A(n6288), .B(n3737), .Z(n6390) );
  CND2X1 U7496 ( .A(n6290), .B(n3731), .Z(n6392) );
  CND2X1 U7497 ( .A(n4572), .B(n3190), .Z(n4623) );
  CND2X1 U7498 ( .A(n5666), .B(n3194), .Z(n5684) );
  CND2X1 U7499 ( .A(n4526), .B(n4224), .Z(n4569) );
  CND2X1 U7500 ( .A(n4509), .B(n4225), .Z(n4532) );
  CND2X1 U7501 ( .A(n5693), .B(n4222), .Z(n5734) );
  CND2X1 U7502 ( .A(n4507), .B(n4225), .Z(n4531) );
  CND2X1 U7503 ( .A(n4464), .B(n3188), .Z(n4496) );
  CND2X1 U7504 ( .A(n4678), .B(n4224), .Z(n4714) );
  CND2X1 U7505 ( .A(n4524), .B(n4224), .Z(n4568) );
  CND2X1 U7506 ( .A(n5714), .B(n4221), .Z(n5749) );
  CND2X1 U7507 ( .A(n5702), .B(n4221), .Z(n5740) );
  CND2X1 U7508 ( .A(n5696), .B(n4221), .Z(n5736) );
  CND2X1 U7509 ( .A(n5151), .B(n4222), .Z(n5185) );
  CND2X1 U7510 ( .A(n5148), .B(n4222), .Z(n5183) );
  CND2X1 U7511 ( .A(n5138), .B(n4222), .Z(n5177) );
  CND2X1 U7512 ( .A(n5135), .B(n4222), .Z(n5175) );
  CND2X1 U7513 ( .A(n5132), .B(n4223), .Z(n5173) );
  CND2X1 U7514 ( .A(n4662), .B(n4223), .Z(n4734) );
  CND2X1 U7515 ( .A(n4648), .B(n4223), .Z(n4726) );
  CND2X1 U7516 ( .A(n4684), .B(n4223), .Z(n4718) );
  CND2X1 U7517 ( .A(n4530), .B(n4224), .Z(n4571) );
  CND2X1 U7518 ( .A(n4656), .B(n4223), .Z(n4730) );
  CND2X1 U7519 ( .A(n4645), .B(n3893), .Z(n4689) );
  CND2X1 U7520 ( .A(n5532), .B(n3892), .Z(n5588) );
  CND2X1 U7521 ( .A(n6094), .B(n3891), .Z(n6126) );
  CND2X1 U7522 ( .A(n6092), .B(n3895), .Z(n6123) );
  CND2X1 U7523 ( .A(n6088), .B(n3892), .Z(n6119) );
  CND2X1 U7524 ( .A(n6083), .B(n3895), .Z(n6115) );
  CND2X1 U7525 ( .A(n6079), .B(n3894), .Z(n6111) );
  CND2X1 U7526 ( .A(n6075), .B(n3894), .Z(n6107) );
  CND2X1 U7527 ( .A(n6070), .B(n3893), .Z(n6103) );
  CND2X1 U7528 ( .A(n6065), .B(n3891), .Z(n6099) );
  CND2X1 U7529 ( .A(n5544), .B(n3893), .Z(n5602) );
  CND2X1 U7530 ( .A(n5538), .B(n3892), .Z(n5595) );
  CND2X1 U7531 ( .A(n5526), .B(n3891), .Z(n5581) );
  CND2X1 U7532 ( .A(n5514), .B(n3891), .Z(n5565) );
  CND2X1 U7533 ( .A(n5508), .B(n3895), .Z(n5558) );
  CND2X1 U7534 ( .A(n5501), .B(n3895), .Z(n5551) );
  CND2X1 U7535 ( .A(n4982), .B(n3894), .Z(n5038) );
  CND2X1 U7536 ( .A(n4963), .B(n3893), .Z(n5017) );
  CND2X1 U7537 ( .A(n4957), .B(n3893), .Z(n5010) );
  CND2X1 U7538 ( .A(n4939), .B(n3892), .Z(n4989) );
  CND2X1 U7539 ( .A(n4687), .B(n3891), .Z(n4747) );
  CND2X1 U7540 ( .A(n4681), .B(n3891), .Z(n4744) );
  CND2X1 U7541 ( .A(n4675), .B(n3895), .Z(n4739) );
  CND2X1 U7542 ( .A(n5520), .B(n3895), .Z(n5574) );
  CIVX2 U7543 ( .A(n4299), .Z(n4268) );
  CIVX2 U7544 ( .A(n4299), .Z(n4269) );
  CND2X1 U7545 ( .A(n4520), .B(n4225), .Z(n4533) );
  CND2X1 U7546 ( .A(n5129), .B(n4223), .Z(n5171) );
  CND2X1 U7547 ( .A(n4522), .B(n4225), .Z(n4534) );
  CND2X1 U7548 ( .A(n4528), .B(n4224), .Z(n4570) );
  CND2X1 U7549 ( .A(n6291), .B(n3724), .Z(n6391) );
  CND2X1 U7550 ( .A(n6286), .B(n3730), .Z(n6387) );
  CND2X1 U7551 ( .A(n6284), .B(n3730), .Z(n6385) );
  CND2X1 U7552 ( .A(n6282), .B(n3729), .Z(n6383) );
  CND2X1 U7553 ( .A(n6280), .B(n3723), .Z(n6381) );
  CND2X1 U7554 ( .A(n6278), .B(n3723), .Z(n6378) );
  CND2X1 U7555 ( .A(n6276), .B(n3728), .Z(n6376) );
  CND2X1 U7556 ( .A(n6265), .B(n3728), .Z(n6366) );
  CND2X1 U7557 ( .A(n6263), .B(n3727), .Z(n6364) );
  CND2X1 U7558 ( .A(n6289), .B(n3724), .Z(n6389) );
  CND2X1 U7559 ( .A(n6270), .B(n3723), .Z(n6370) );
  CND2X1 U7560 ( .A(n6274), .B(n3729), .Z(n6374) );
  CND2X1 U7561 ( .A(n6272), .B(n3728), .Z(n6372) );
  CND2X1 U7562 ( .A(n4826), .B(n3736), .Z(n4946) );
  CND2X1 U7563 ( .A(n4823), .B(n3737), .Z(n4940) );
  CND2X1 U7564 ( .A(n4815), .B(n3733), .Z(n4921) );
  CND2X1 U7565 ( .A(n6257), .B(n3726), .Z(n6357) );
  CND2X1 U7566 ( .A(n6268), .B(n3725), .Z(n6368) );
  CND2X1 U7567 ( .A(n6255), .B(n3726), .Z(n6355) );
  CND2X1 U7568 ( .A(n4842), .B(n3733), .Z(n4997) );
  CND2X1 U7569 ( .A(n4836), .B(n3739), .Z(n4976) );
  CND2X1 U7570 ( .A(n4834), .B(n3737), .Z(n4970) );
  CND2X1 U7571 ( .A(n4830), .B(n3737), .Z(n4958) );
  CND2X1 U7572 ( .A(n4828), .B(n3731), .Z(n4952) );
  CND2X1 U7573 ( .A(n6261), .B(n3722), .Z(n6362) );
  CND2X1 U7574 ( .A(n6259), .B(n3728), .Z(n6360) );
  CND2X1 U7575 ( .A(n6253), .B(n3726), .Z(n6353) );
  CND2X1 U7576 ( .A(n6251), .B(n3727), .Z(n6351) );
  CND2X1 U7577 ( .A(n6249), .B(n3726), .Z(n6349) );
  CND2X1 U7578 ( .A(n6247), .B(n3728), .Z(n6347) );
  CND2X1 U7579 ( .A(n6244), .B(n3721), .Z(n6345) );
  CND2X1 U7580 ( .A(n6242), .B(n3727), .Z(n6343) );
  CND2X1 U7581 ( .A(n4870), .B(n3731), .Z(n5089) );
  CND2X1 U7582 ( .A(n4868), .B(n3736), .Z(n5082) );
  CND2X1 U7583 ( .A(n4865), .B(n3736), .Z(n5075) );
  CND2X1 U7584 ( .A(n4863), .B(n3731), .Z(n5068) );
  CND2X1 U7585 ( .A(n4861), .B(n3739), .Z(n5061) );
  CND2X1 U7586 ( .A(n4859), .B(n3732), .Z(n5054) );
  CND2X1 U7587 ( .A(n4857), .B(n3738), .Z(n5046) );
  CND2X1 U7588 ( .A(n4855), .B(n3734), .Z(n5039) );
  CND2X1 U7589 ( .A(n4853), .B(n3731), .Z(n5032) );
  CND2X1 U7590 ( .A(n4851), .B(n3740), .Z(n5025) );
  CND2X1 U7591 ( .A(n4849), .B(n3732), .Z(n5018) );
  CND2X1 U7592 ( .A(n4847), .B(n3738), .Z(n5011) );
  CND2X1 U7593 ( .A(n4844), .B(n3737), .Z(n5004) );
  CND2X1 U7594 ( .A(n4840), .B(n3735), .Z(n4990) );
  CND2X1 U7595 ( .A(n4838), .B(n3733), .Z(n4983) );
  CND2X1 U7596 ( .A(n5741), .B(n3207), .Z(n5808) );
  CND2X1 U7597 ( .A(n5739), .B(n3205), .Z(n5806) );
  CND2X1 U7598 ( .A(n5707), .B(n3203), .Z(n5776) );
  CND2X1 U7599 ( .A(n12699), .B(n4010), .Z(n12709) );
  CND2X1 U7600 ( .A(n9627), .B(n4010), .Z(n9637) );
  CND2X1 U7601 ( .A(n12702), .B(n4010), .Z(n12711) );
  CND2X1 U7602 ( .A(n5711), .B(n4221), .Z(n5747) );
  CANR2X1 U7603 ( .A(N3106), .B(n3592), .C(N2072), .D(n3637), .Z(n2112) );
  CND2X1 U7604 ( .A(n2110), .B(n2111), .Z(N10355) );
  CANR2X1 U7605 ( .A(N6226), .B(n3592), .C(n3760), .D(n3637), .Z(n2116) );
  CND2X1 U7606 ( .A(n2108), .B(n2109), .Z(N10356) );
  CANR2X1 U7607 ( .A(N6225), .B(n3592), .C(n3892), .D(n3637), .Z(n2118) );
  CNIVX1 U7608 ( .A(n4006), .Z(n4180) );
  CNIVX1 U7609 ( .A(n4006), .Z(n4179) );
  CNIVX1 U7610 ( .A(n4006), .Z(n4181) );
  CNIVX1 U7611 ( .A(n4006), .Z(n4183) );
  CNIVX1 U7612 ( .A(n4007), .Z(n4187) );
  CNIVX1 U7613 ( .A(n4007), .Z(n4188) );
  CNIVX1 U7614 ( .A(n4005), .Z(n4175) );
  CNIVX1 U7615 ( .A(n4005), .Z(n4173) );
  CNIVX1 U7616 ( .A(n4005), .Z(n4174) );
  CNIVX1 U7617 ( .A(n4005), .Z(n4176) );
  CNIVX1 U7618 ( .A(n4006), .Z(n4182) );
  CNIVX1 U7619 ( .A(n4006), .Z(n4184) );
  CNIVX1 U7620 ( .A(n4007), .Z(n4186) );
  CNIVX1 U7621 ( .A(n4007), .Z(n4189) );
  CNIVX1 U7622 ( .A(n4009), .Z(n4201) );
  CNIVX1 U7623 ( .A(n3991), .Z(n4073) );
  CNIVX1 U7624 ( .A(n4000), .Z(n4137) );
  CNIVX1 U7625 ( .A(n3982), .Z(n4011) );
  CNIVX1 U7626 ( .A(n3991), .Z(n4075) );
  CNIVX1 U7627 ( .A(n4000), .Z(n4139) );
  CNIVX1 U7628 ( .A(n3982), .Z(n4012) );
  CNIVX1 U7629 ( .A(n3991), .Z(n4076) );
  CNIVX1 U7630 ( .A(n4000), .Z(n4140) );
  CNIVX1 U7631 ( .A(n3982), .Z(n4013) );
  CNIVX1 U7632 ( .A(n3991), .Z(n4077) );
  CNIVX1 U7633 ( .A(n4000), .Z(n4141) );
  CNIVX1 U7634 ( .A(n3982), .Z(n4014) );
  CNIVX1 U7635 ( .A(n3991), .Z(n4078) );
  CNIVX1 U7636 ( .A(n4000), .Z(n4142) );
  CNIVX1 U7637 ( .A(n3982), .Z(n4015) );
  CNIVX1 U7638 ( .A(n3991), .Z(n4079) );
  CNIVX1 U7639 ( .A(n4001), .Z(n4143) );
  CNIVX1 U7640 ( .A(n3982), .Z(n4016) );
  CNIVX1 U7641 ( .A(n3992), .Z(n4080) );
  CNIVX1 U7642 ( .A(n4001), .Z(n4144) );
  CNIVX1 U7643 ( .A(n4009), .Z(n4200) );
  CNIVX1 U7644 ( .A(n4000), .Z(n4136) );
  CNIVX1 U7645 ( .A(n3990), .Z(n4072) );
  CNIVX1 U7646 ( .A(n4001), .Z(n4145) );
  CNIVX1 U7647 ( .A(n3992), .Z(n4081) );
  CNIVX1 U7648 ( .A(n3983), .Z(n4017) );
  CNIVX1 U7649 ( .A(n4001), .Z(n4146) );
  CNIVX1 U7650 ( .A(n3992), .Z(n4082) );
  CNIVX1 U7651 ( .A(n3983), .Z(n4018) );
  CNIVX1 U7652 ( .A(n3983), .Z(n4019) );
  CNIVX1 U7653 ( .A(n4001), .Z(n4147) );
  CNIVX1 U7654 ( .A(n3992), .Z(n4083) );
  CNIVX1 U7655 ( .A(n4001), .Z(n4148) );
  CNIVX1 U7656 ( .A(n3992), .Z(n4084) );
  CNIVX1 U7657 ( .A(n3983), .Z(n4020) );
  CNIVX1 U7658 ( .A(n3983), .Z(n4021) );
  CNIVX1 U7659 ( .A(n4001), .Z(n4149) );
  CNIVX1 U7660 ( .A(n3992), .Z(n4085) );
  CNIVX1 U7661 ( .A(n4002), .Z(n4150) );
  CNIVX1 U7662 ( .A(n3992), .Z(n4086) );
  CNIVX1 U7663 ( .A(n3983), .Z(n4022) );
  CNIVX1 U7664 ( .A(n3993), .Z(n4087) );
  CNIVX1 U7665 ( .A(n3983), .Z(n4023) );
  CNIVX1 U7666 ( .A(n4002), .Z(n4151) );
  CNIVX1 U7667 ( .A(n4002), .Z(n4152) );
  CNIVX1 U7668 ( .A(n3993), .Z(n4088) );
  CNIVX1 U7669 ( .A(n3984), .Z(n4024) );
  CNIVX1 U7670 ( .A(n3993), .Z(n4089) );
  CNIVX1 U7671 ( .A(n3984), .Z(n4025) );
  CNIVX1 U7672 ( .A(n4002), .Z(n4153) );
  CNIVX1 U7673 ( .A(n4002), .Z(n4154) );
  CNIVX1 U7674 ( .A(n3993), .Z(n4090) );
  CNIVX1 U7675 ( .A(n3984), .Z(n4026) );
  CNIVX1 U7676 ( .A(n4002), .Z(n4155) );
  CNIVX1 U7677 ( .A(n3993), .Z(n4091) );
  CNIVX1 U7678 ( .A(n3984), .Z(n4027) );
  CNIVX1 U7679 ( .A(n4002), .Z(n4156) );
  CNIVX1 U7680 ( .A(n3993), .Z(n4092) );
  CNIVX1 U7681 ( .A(n3984), .Z(n4028) );
  CNIVX1 U7682 ( .A(n4003), .Z(n4157) );
  CNIVX1 U7683 ( .A(n3993), .Z(n4093) );
  CNIVX1 U7684 ( .A(n3984), .Z(n4029) );
  CNIVX1 U7685 ( .A(n3984), .Z(n4030) );
  CNIVX1 U7686 ( .A(n4003), .Z(n4158) );
  CNIVX1 U7687 ( .A(n3994), .Z(n4094) );
  CNIVX1 U7688 ( .A(n4003), .Z(n4160) );
  CNIVX1 U7689 ( .A(n3994), .Z(n4096) );
  CNIVX1 U7690 ( .A(n4003), .Z(n4161) );
  CNIVX1 U7691 ( .A(n3994), .Z(n4097) );
  CNIVX1 U7692 ( .A(n3985), .Z(n4033) );
  CNIVX1 U7693 ( .A(n3994), .Z(n4098) );
  CNIVX1 U7694 ( .A(n3985), .Z(n4034) );
  CNIVX1 U7695 ( .A(n4003), .Z(n4162) );
  CNIVX1 U7696 ( .A(n4003), .Z(n4163) );
  CNIVX1 U7697 ( .A(n3994), .Z(n4099) );
  CNIVX1 U7698 ( .A(n3985), .Z(n4035) );
  CNIVX1 U7699 ( .A(n3994), .Z(n4100) );
  CNIVX1 U7700 ( .A(n3985), .Z(n4036) );
  CNIVX1 U7701 ( .A(n4004), .Z(n4164) );
  CNIVX1 U7702 ( .A(n4004), .Z(n4165) );
  CNIVX1 U7703 ( .A(n3995), .Z(n4101) );
  CNIVX1 U7704 ( .A(n3985), .Z(n4037) );
  CNIVX1 U7705 ( .A(n4004), .Z(n4166) );
  CNIVX1 U7706 ( .A(n3995), .Z(n4102) );
  CNIVX1 U7707 ( .A(n3986), .Z(n4038) );
  CNIVX1 U7708 ( .A(n4004), .Z(n4167) );
  CNIVX1 U7709 ( .A(n3995), .Z(n4103) );
  CNIVX1 U7710 ( .A(n3986), .Z(n4039) );
  CNIVX1 U7711 ( .A(n4004), .Z(n4168) );
  CNIVX1 U7712 ( .A(n3995), .Z(n4104) );
  CNIVX1 U7713 ( .A(n3986), .Z(n4040) );
  CNIVX1 U7714 ( .A(n3986), .Z(n4041) );
  CNIVX1 U7715 ( .A(n4004), .Z(n4169) );
  CNIVX1 U7716 ( .A(n3995), .Z(n4105) );
  CNIVX1 U7717 ( .A(n4004), .Z(n4170) );
  CNIVX1 U7718 ( .A(n3995), .Z(n4106) );
  CNIVX1 U7719 ( .A(n3986), .Z(n4042) );
  CNIVX1 U7720 ( .A(n3986), .Z(n4043) );
  CNIVX1 U7721 ( .A(n4005), .Z(n4171) );
  CNIVX1 U7722 ( .A(n3995), .Z(n4107) );
  CNIVX1 U7723 ( .A(n3996), .Z(n4108) );
  CNIVX1 U7724 ( .A(n3986), .Z(n4044) );
  CNIVX1 U7725 ( .A(n3996), .Z(n4109) );
  CNIVX1 U7726 ( .A(n3987), .Z(n4045) );
  CNIVX1 U7727 ( .A(n3996), .Z(n4110) );
  CNIVX1 U7728 ( .A(n3987), .Z(n4046) );
  CNIVX1 U7729 ( .A(n3996), .Z(n4111) );
  CNIVX1 U7730 ( .A(n3987), .Z(n4047) );
  CNIVX1 U7731 ( .A(n3996), .Z(n4112) );
  CNIVX1 U7732 ( .A(n3987), .Z(n4048) );
  CNIVX1 U7733 ( .A(n3996), .Z(n4113) );
  CNIVX1 U7734 ( .A(n3987), .Z(n4049) );
  CNIVX1 U7735 ( .A(n3997), .Z(n4115) );
  CNIVX1 U7736 ( .A(n3987), .Z(n4051) );
  CNIVX1 U7737 ( .A(n3997), .Z(n4116) );
  CNIVX1 U7738 ( .A(n3988), .Z(n4052) );
  CNIVX1 U7739 ( .A(n3997), .Z(n4117) );
  CNIVX1 U7740 ( .A(n3988), .Z(n4053) );
  CNIVX1 U7741 ( .A(n3997), .Z(n4118) );
  CNIVX1 U7742 ( .A(n3988), .Z(n4054) );
  CNIVX1 U7743 ( .A(n3997), .Z(n4119) );
  CNIVX1 U7744 ( .A(n3988), .Z(n4055) );
  CNIVX1 U7745 ( .A(n3997), .Z(n4120) );
  CNIVX1 U7746 ( .A(n3988), .Z(n4056) );
  CNIVX1 U7747 ( .A(n3998), .Z(n4122) );
  CNIVX1 U7748 ( .A(n3988), .Z(n4058) );
  CNIVX1 U7749 ( .A(n3998), .Z(n4123) );
  CNIVX1 U7750 ( .A(n3989), .Z(n4059) );
  CNIVX1 U7751 ( .A(n3998), .Z(n4124) );
  CNIVX1 U7752 ( .A(n3989), .Z(n4060) );
  CNIVX1 U7753 ( .A(n3998), .Z(n4125) );
  CNIVX1 U7754 ( .A(n3989), .Z(n4061) );
  CNIVX1 U7755 ( .A(n4007), .Z(n4190) );
  CNIVX1 U7756 ( .A(n3998), .Z(n4126) );
  CNIVX1 U7757 ( .A(n3989), .Z(n4062) );
  CNIVX1 U7758 ( .A(n4007), .Z(n4191) );
  CNIVX1 U7759 ( .A(n3998), .Z(n4127) );
  CNIVX1 U7760 ( .A(n3989), .Z(n4063) );
  CNIVX1 U7761 ( .A(n3999), .Z(n4129) );
  CNIVX1 U7762 ( .A(n3989), .Z(n4065) );
  CNIVX1 U7763 ( .A(n3999), .Z(n4130) );
  CNIVX1 U7764 ( .A(n3990), .Z(n4066) );
  CNIVX1 U7765 ( .A(n4008), .Z(n4194) );
  CNIVX1 U7766 ( .A(n4008), .Z(n4195) );
  CNIVX1 U7767 ( .A(n3999), .Z(n4131) );
  CNIVX1 U7768 ( .A(n3990), .Z(n4067) );
  CNIVX1 U7769 ( .A(n4008), .Z(n4197) );
  CNIVX1 U7770 ( .A(n3999), .Z(n4133) );
  CNIVX1 U7771 ( .A(n3990), .Z(n4069) );
  CNIVX1 U7772 ( .A(n4006), .Z(n4178) );
  CNIVX1 U7773 ( .A(n3999), .Z(n4134) );
  CNIVX1 U7774 ( .A(n3996), .Z(n4114) );
  CNIVX1 U7775 ( .A(n3990), .Z(n4070) );
  CNIVX1 U7776 ( .A(n3987), .Z(n4050) );
  CNIVX1 U7777 ( .A(n3999), .Z(n4135) );
  CNIVX1 U7778 ( .A(n3997), .Z(n4121) );
  CNIVX1 U7779 ( .A(n3990), .Z(n4071) );
  CNIVX1 U7780 ( .A(n3988), .Z(n4057) );
  CNIVX1 U7781 ( .A(n4008), .Z(n4196) );
  CNIVX1 U7782 ( .A(n4008), .Z(n4192) );
  CNIVX1 U7783 ( .A(n3999), .Z(n4132) );
  CNIVX1 U7784 ( .A(n3998), .Z(n4128) );
  CNIVX1 U7785 ( .A(n3990), .Z(n4068) );
  CNIVX1 U7786 ( .A(n3989), .Z(n4064) );
  CNIVX1 U7787 ( .A(n4000), .Z(n4138) );
  CNIVX1 U7788 ( .A(n3991), .Z(n4074) );
  CNIVX1 U7789 ( .A(n4003), .Z(n4159) );
  CNIVX1 U7790 ( .A(n3994), .Z(n4095) );
  CNIVX1 U7791 ( .A(n3985), .Z(n4032) );
  CNIVX1 U7792 ( .A(n3985), .Z(n4031) );
  CNIVX1 U7793 ( .A(n3982), .Z(n4010) );
  CNIVX1 U7794 ( .A(n4009), .Z(n4199) );
  CNIVX1 U7795 ( .A(n4005), .Z(n4172) );
  CNIVX1 U7796 ( .A(n4005), .Z(n4177) );
  CNIVX1 U7797 ( .A(n4007), .Z(n4185) );
  CIVX2 U7798 ( .A(n4300), .Z(n4288) );
  CIVX2 U7799 ( .A(n4300), .Z(n4287) );
  CIVX2 U7800 ( .A(n4300), .Z(n4290) );
  CIVX2 U7801 ( .A(n4300), .Z(n4291) );
  CIVX2 U7802 ( .A(n4300), .Z(n4292) );
  CIVX2 U7803 ( .A(n4298), .Z(n4262) );
  CIVX2 U7804 ( .A(n4298), .Z(n4263) );
  CIVX2 U7805 ( .A(n4298), .Z(n4264) );
  CIVX2 U7806 ( .A(n4298), .Z(n4265) );
  CIVX2 U7807 ( .A(n4298), .Z(n4266) );
  CIVX2 U7808 ( .A(n4299), .Z(n4271) );
  CIVX2 U7809 ( .A(n4299), .Z(n4273) );
  CIVX2 U7810 ( .A(n4299), .Z(n4274) );
  CIVX2 U7811 ( .A(n4299), .Z(n4275) );
  CIVX2 U7812 ( .A(n4299), .Z(n4276) );
  CIVX2 U7813 ( .A(n4299), .Z(n4277) );
  CIVX2 U7814 ( .A(n4299), .Z(n4278) );
  CIVX2 U7815 ( .A(n4296), .Z(n4247) );
  CIVX2 U7816 ( .A(n4297), .Z(n4250) );
  CIVX2 U7817 ( .A(n4299), .Z(n4279) );
  CIVX2 U7818 ( .A(n4300), .Z(n4283) );
  CIVX2 U7819 ( .A(n4300), .Z(n4289) );
  CIVX2 U7820 ( .A(n4379), .Z(n4366) );
  CIVX2 U7821 ( .A(n4379), .Z(n4367) );
  CIVX2 U7822 ( .A(n4382), .Z(n4339) );
  CIVX2 U7823 ( .A(n4382), .Z(n4340) );
  CIVX2 U7824 ( .A(n4381), .Z(n4342) );
  CIVX2 U7825 ( .A(n4381), .Z(n4343) );
  CIVX2 U7826 ( .A(n4381), .Z(n4344) );
  CIVX2 U7827 ( .A(n4381), .Z(n4346) );
  CIVX2 U7828 ( .A(n4381), .Z(n4347) );
  CIVX2 U7829 ( .A(n4384), .Z(n4308) );
  CIVX2 U7830 ( .A(n4381), .Z(n4348) );
  CIVX2 U7831 ( .A(n4384), .Z(n4309) );
  CIVX2 U7832 ( .A(n4381), .Z(n4349) );
  CIVX2 U7833 ( .A(n4384), .Z(n4310) );
  CIVX2 U7834 ( .A(n4381), .Z(n4350) );
  CIVX2 U7835 ( .A(n4384), .Z(n4311) );
  CIVX2 U7836 ( .A(n4381), .Z(n4351) );
  CIVX2 U7837 ( .A(n4384), .Z(n4312) );
  CIVX2 U7838 ( .A(n4384), .Z(n4313) );
  CIVX2 U7839 ( .A(n4383), .Z(n4322) );
  CIVX2 U7840 ( .A(n4384), .Z(n4314) );
  CIVX2 U7841 ( .A(n4383), .Z(n4323) );
  CIVX2 U7842 ( .A(n4384), .Z(n4315) );
  CIVX2 U7843 ( .A(n4383), .Z(n4324) );
  CIVX2 U7844 ( .A(n4384), .Z(n4316) );
  CIVX2 U7845 ( .A(n4383), .Z(n4325) );
  CIVX2 U7846 ( .A(n4384), .Z(n4317) );
  CIVX2 U7847 ( .A(n4383), .Z(n4326) );
  CIVX2 U7848 ( .A(n4384), .Z(n4318) );
  CIVX2 U7849 ( .A(n4383), .Z(n4327) );
  CIVX2 U7850 ( .A(n4383), .Z(n4328) );
  CIVX2 U7851 ( .A(n4383), .Z(n4319) );
  CIVX2 U7852 ( .A(n4382), .Z(n4331) );
  CIVX2 U7853 ( .A(n4383), .Z(n4320) );
  CIVX2 U7854 ( .A(n4382), .Z(n4332) );
  CIVX2 U7855 ( .A(n4383), .Z(n4321) );
  CIVX2 U7856 ( .A(n4382), .Z(n4333) );
  CIVX2 U7857 ( .A(n4382), .Z(n4334) );
  CIVX2 U7858 ( .A(n4382), .Z(n4335) );
  CIVX2 U7859 ( .A(n4382), .Z(n4336) );
  CIVX2 U7860 ( .A(n4382), .Z(n4337) );
  CIVX2 U7861 ( .A(n4382), .Z(n4338) );
  CIVX2 U7862 ( .A(n4379), .Z(n4369) );
  CIVX2 U7863 ( .A(n4379), .Z(n4370) );
  CIVX2 U7864 ( .A(n4379), .Z(n4371) );
  CIVX2 U7865 ( .A(n4379), .Z(n4372) );
  CIVX2 U7866 ( .A(n4379), .Z(n4373) );
  CIVX2 U7867 ( .A(n4379), .Z(n4374) );
  CIVX2 U7868 ( .A(n4379), .Z(n4375) );
  CIVX2 U7869 ( .A(n4380), .Z(n4354) );
  CIVX2 U7870 ( .A(n4380), .Z(n4355) );
  CIVX2 U7871 ( .A(n4380), .Z(n4356) );
  CIVX2 U7872 ( .A(n4380), .Z(n4358) );
  CIVX2 U7873 ( .A(n4380), .Z(n4363) );
  CIVX2 U7874 ( .A(n4380), .Z(n4359) );
  CIVX2 U7875 ( .A(n4380), .Z(n4360) );
  CIVX2 U7876 ( .A(n4380), .Z(n4361) );
  CIVX2 U7877 ( .A(n4380), .Z(n4362) );
  CIVX2 U7878 ( .A(n4380), .Z(n4364) );
  CIVX2 U7879 ( .A(n4379), .Z(n4365) );
  CIVX2 U7880 ( .A(n4380), .Z(n4357) );
  CIVX2 U7881 ( .A(n4379), .Z(n4368) );
  CIVX2 U7882 ( .A(n4381), .Z(n4345) );
  CIVX2 U7883 ( .A(n4297), .Z(n4251) );
  CIVX2 U7884 ( .A(n4296), .Z(n4241) );
  CIVX2 U7885 ( .A(n4296), .Z(n4246) );
  CIVX2 U7886 ( .A(n4299), .Z(n4280) );
  CIVX2 U7887 ( .A(n4300), .Z(n4284) );
  CIVX2 U7888 ( .A(n4297), .Z(n4252) );
  CIVX2 U7889 ( .A(n4297), .Z(n4253) );
  CIVX2 U7890 ( .A(n4298), .Z(n4261) );
  CIVX2 U7891 ( .A(n4297), .Z(n4254) );
  CIVX2 U7892 ( .A(n4297), .Z(n4255) );
  CIVX2 U7893 ( .A(n4298), .Z(n4258) );
  CIVX2 U7894 ( .A(n4298), .Z(n4259) );
  CIVX2 U7895 ( .A(n4300), .Z(n4285) );
  CIVX2 U7896 ( .A(n4296), .Z(n4242) );
  CNIVX1 U7897 ( .A(n4009), .Z(n4202) );
  CIVX2 U7898 ( .A(n4300), .Z(n4286) );
  CIVX2 U7899 ( .A(n4296), .Z(n4244) );
  CIVX2 U7900 ( .A(n4296), .Z(n4245) );
  CIVX2 U7901 ( .A(n4297), .Z(n4248) );
  CIVX2 U7902 ( .A(n4300), .Z(n4281) );
  CIVX2 U7903 ( .A(n4300), .Z(n4282) );
  CIVX2 U7904 ( .A(n4380), .Z(n4353) );
  CIVX2 U7905 ( .A(n4381), .Z(n4341) );
  CIVX2 U7906 ( .A(n4380), .Z(n4352) );
  CIVX2 U7907 ( .A(n4382), .Z(n4329) );
  CIVX2 U7908 ( .A(n4382), .Z(n4330) );
  CIVX2 U7909 ( .A(n4384), .Z(n4307) );
  CIVX2 U7910 ( .A(n4296), .Z(n4239) );
  CIVX2 U7911 ( .A(n4297), .Z(n4249) );
  CIVX2 U7912 ( .A(n4298), .Z(n4260) );
  CIVX2 U7913 ( .A(n4296), .Z(n4240) );
  CIVX2 U7914 ( .A(n4296), .Z(n4243) );
  CIVX2 U7915 ( .A(n4298), .Z(n4257) );
  CIVX2 U7916 ( .A(n4298), .Z(n4256) );
  CNIVX1 U7917 ( .A(n3755), .Z(n3762) );
  CNIVXL U7918 ( .A(n3248), .Z(n3648) );
  CNIVXL U7919 ( .A(n3249), .Z(n3649) );
  CNIVXL U7920 ( .A(n3248), .Z(n3650) );
  CNIVXL U7921 ( .A(n3249), .Z(n3651) );
  CNIVXL U7922 ( .A(n3248), .Z(n3647) );
  CNIVXL U7923 ( .A(n3249), .Z(n3646) );
  CNIVXL U7924 ( .A(n3248), .Z(n3645) );
  CNIVXL U7925 ( .A(n3249), .Z(n3675) );
  CNIVXL U7926 ( .A(n3248), .Z(n3676) );
  CNIVX1 U7927 ( .A(n3248), .Z(n3679) );
  CNIVX1 U7928 ( .A(n3249), .Z(n3678) );
  CNIVX1 U7929 ( .A(n3249), .Z(n3681) );
  CNIVX1 U7930 ( .A(n3248), .Z(n3680) );
  CENX1 U7931 ( .A(n4400), .B(n3267), .Z(N3109) );
  CENX1 U7932 ( .A(N431), .B(n3743), .Z(n3714) );
  CNIVX1 U7933 ( .A(n3752), .Z(n3891) );
  CMXI2X1 U7934 ( .A0(N8272), .A1(N8271), .S(n3859), .Z(n13737) );
  CMXI2X1 U7935 ( .A0(N8274), .A1(N8273), .S(n3859), .Z(n13740) );
  CMXI2X1 U7936 ( .A0(N8273), .A1(N8272), .S(n3857), .Z(n13400) );
  CMXI2X1 U7937 ( .A0(N8275), .A1(N8274), .S(n3857), .Z(n13403) );
  CMX2X1 U7938 ( .A0(n3268), .A1(n3269), .S(n4175), .Z(n13864) );
  CMXI2X1 U7939 ( .A0(N7832), .A1(N7831), .S(n3862), .Z(n3268) );
  CMXI2X1 U7940 ( .A0(N7834), .A1(N7833), .S(n3871), .Z(n3269) );
  CNIVX1 U7941 ( .A(n3754), .Z(n3892) );
  CNIVX1 U7942 ( .A(n3754), .Z(n3893) );
  CNR2X1 U7943 ( .A(n4620), .B(n3247), .Z(n4675) );
  CNR2X1 U7944 ( .A(n4491), .B(n3896), .Z(n4526) );
  CNR2X1 U7945 ( .A(n5676), .B(n3896), .Z(n5705) );
  CNR2X1 U7946 ( .A(n4486), .B(n3896), .Z(n4524) );
  CNR2X1 U7947 ( .A(n5688), .B(n3896), .Z(n5714) );
  CNR2X1 U7948 ( .A(n5684), .B(n3896), .Z(n5711) );
  CNR2X1 U7949 ( .A(n5680), .B(n3896), .Z(n5708) );
  CNR2X1 U7950 ( .A(n5125), .B(n3896), .Z(n5151) );
  CNR2X1 U7951 ( .A(n5121), .B(n3896), .Z(n5148) );
  CNR2X1 U7952 ( .A(n4633), .B(n3896), .Z(n4662) );
  CNR2X1 U7953 ( .A(n4496), .B(n3896), .Z(n4528) );
  CNR2X1 U7954 ( .A(n4501), .B(n3896), .Z(n4530) );
  CNR2X1 U7955 ( .A(n4623), .B(n3896), .Z(n4656) );
  CNR2X1 U7956 ( .A(n6049), .B(n4219), .Z(n6070) );
  CNR2X1 U7957 ( .A(n4925), .B(n4219), .Z(n4945) );
  CNR2X1 U7958 ( .A(n5485), .B(n4217), .Z(n5508) );
  CNR2X1 U7959 ( .A(n4630), .B(n3246), .Z(n4681) );
  CNR2IX1 U7960 ( .B(n6217), .A(n3200), .Z(n6284) );
  CNR2IX1 U7961 ( .B(n4771), .A(n3216), .Z(n4837) );
  CNIVX1 U7962 ( .A(n3753), .Z(n3895) );
  CNIVX1 U7963 ( .A(n4436), .Z(n4207) );
  CNIVX1 U7964 ( .A(n3753), .Z(n3894) );
  CND2X1 U7965 ( .A(n3722), .B(n5823), .Z(n5925) );
  CND2X1 U7966 ( .A(n5823), .B(n3734), .Z(n5996) );
  CND2X1 U7967 ( .A(n3728), .B(n5275), .Z(n5378) );
  CND2X1 U7968 ( .A(n5275), .B(n3736), .Z(n5448) );
  CIVX2 U7969 ( .A(n3754), .Z(n4226) );
  CNIVX1 U7970 ( .A(n4436), .Z(n4203) );
  CNIVX1 U7971 ( .A(n4436), .Z(n4209) );
  CNIVX1 U7972 ( .A(n4436), .Z(n4204) );
  CNIVX1 U7973 ( .A(n4436), .Z(n4210) );
  CNIVX1 U7974 ( .A(n4436), .Z(n4205) );
  CNIVX1 U7975 ( .A(n4436), .Z(n4208) );
  CNIVX1 U7976 ( .A(n4436), .Z(n4206) );
  CND2X1 U7977 ( .A(n6273), .B(n3739), .Z(n6375) );
  CND2X1 U7978 ( .A(n5090), .B(n4407), .Z(n4441) );
  CND2X1 U7979 ( .A(n5654), .B(n4410), .Z(n5660) );
  CND2X1 U7980 ( .A(n6027), .B(n4408), .Z(n6030) );
  CND2X1 U7981 ( .A(n5464), .B(n4410), .Z(n5467) );
  CNR2IX1 U7982 ( .B(N7256), .A(n3859), .Z(n9630) );
  CND2X1 U7983 ( .A(n5492), .B(n4394), .Z(n4558) );
  CND2X1 U7984 ( .A(n5033), .B(n4398), .Z(n5041) );
  CND2X1 U7985 ( .A(n4947), .B(n4397), .Z(n4954) );
  CND2X1 U7986 ( .A(n5026), .B(n4398), .Z(n5034) );
  CND2X1 U7987 ( .A(n4953), .B(n4397), .Z(n4960) );
  CND2X1 U7988 ( .A(n5504), .B(n4394), .Z(n4556) );
  CND2X1 U7989 ( .A(n5019), .B(n4398), .Z(n5027) );
  CND2X1 U7990 ( .A(n5012), .B(n4398), .Z(n5020) );
  CND2X1 U7991 ( .A(n5473), .B(n4394), .Z(n4562) );
  CND2X1 U7992 ( .A(n5005), .B(n4398), .Z(n5013) );
  CND2X1 U7993 ( .A(n4965), .B(n4397), .Z(n4972) );
  CND2X1 U7994 ( .A(n4998), .B(n4398), .Z(n5006) );
  CND2X1 U7995 ( .A(n5487), .B(n4394), .Z(n4561) );
  CND2X1 U7996 ( .A(n4971), .B(n4397), .Z(n4979) );
  CND2X1 U7997 ( .A(n4978), .B(n4397), .Z(n4985) );
  CND2X1 U7998 ( .A(n5477), .B(n4394), .Z(n4563) );
  CND2X1 U7999 ( .A(n4984), .B(n4397), .Z(n4992) );
  CND2X1 U8000 ( .A(n6029), .B(n4413), .Z(n6033) );
  CND2X1 U8001 ( .A(n5033), .B(n4402), .Z(n4448) );
  CND2X1 U8002 ( .A(n5040), .B(n4402), .Z(n4449) );
  CND2X1 U8003 ( .A(n5026), .B(n4403), .Z(n4451) );
  CND2X1 U8004 ( .A(n4991), .B(n4404), .Z(n4454) );
  CND2X1 U8005 ( .A(n5069), .B(n4401), .Z(n4445) );
  CND2X1 U8006 ( .A(n5062), .B(n4401), .Z(n4444) );
  CND2X1 U8007 ( .A(n5019), .B(n4403), .Z(n4450) );
  CND2X1 U8008 ( .A(n5048), .B(n4402), .Z(n4446) );
  CND2X1 U8009 ( .A(n5012), .B(n4403), .Z(n4453) );
  CND2X1 U8010 ( .A(n5055), .B(n4401), .Z(n4447) );
  CND2X1 U8011 ( .A(n5005), .B(n4404), .Z(n4452) );
  CND2X1 U8012 ( .A(n4998), .B(n4404), .Z(n4455) );
  CND2X1 U8013 ( .A(n4832), .B(n3738), .Z(n4964) );
  CND2X1 U8014 ( .A(n5076), .B(n4411), .Z(n4442) );
  CND2X1 U8015 ( .A(n4984), .B(n4405), .Z(n4457) );
  CND2X1 U8016 ( .A(n4978), .B(n4405), .Z(n4456) );
  CND2X1 U8017 ( .A(n4971), .B(n4405), .Z(n4459) );
  CND2X1 U8018 ( .A(n4965), .B(n4411), .Z(n4458) );
  CND2X1 U8019 ( .A(n4959), .B(n4412), .Z(n4461) );
  CND2X1 U8020 ( .A(n4953), .B(n4407), .Z(n4460) );
  CND2X1 U8021 ( .A(n4947), .B(n4409), .Z(n4463) );
  CND2X1 U8022 ( .A(n4941), .B(n4406), .Z(n4462) );
  CND2X1 U8023 ( .A(n5083), .B(n4412), .Z(n4443) );
  CND2X1 U8024 ( .A(n5625), .B(n4412), .Z(n5633) );
  CND2X1 U8025 ( .A(n5618), .B(n4408), .Z(n5626) );
  CND2X1 U8026 ( .A(n5611), .B(n4410), .Z(n5619) );
  CND2X1 U8027 ( .A(n5583), .B(n4411), .Z(n5591) );
  CND2X1 U8028 ( .A(n5576), .B(n4410), .Z(n5584) );
  CND2X1 U8029 ( .A(n5597), .B(n4411), .Z(n5605) );
  CND2X1 U8030 ( .A(n5590), .B(n4411), .Z(n5598) );
  CND2X1 U8031 ( .A(n5640), .B(n4412), .Z(n5648) );
  CND2X1 U8032 ( .A(n5632), .B(n4412), .Z(n5641) );
  CND2X1 U8033 ( .A(n5647), .B(n4408), .Z(n5655) );
  CND2X1 U8034 ( .A(n5516), .B(n4408), .Z(n5523) );
  CND2X1 U8035 ( .A(n5510), .B(n4408), .Z(n5517) );
  CND2X1 U8036 ( .A(n5504), .B(n4408), .Z(n5511) );
  CND2X1 U8037 ( .A(n5497), .B(n4407), .Z(n5505) );
  CND2X1 U8038 ( .A(n5492), .B(n4407), .Z(n5498) );
  CND2X1 U8039 ( .A(n5487), .B(n4407), .Z(n5493) );
  CND2X1 U8040 ( .A(n5477), .B(n4406), .Z(n5483) );
  CND2X1 U8041 ( .A(n5482), .B(n4406), .Z(n5488) );
  CND2X1 U8042 ( .A(n5569), .B(n4410), .Z(n5577) );
  CND2X1 U8043 ( .A(n5560), .B(n4410), .Z(n5570) );
  CND2X1 U8044 ( .A(n5546), .B(n4409), .Z(n5554) );
  CND2X1 U8045 ( .A(n5553), .B(n4409), .Z(n5561) );
  CND2X1 U8046 ( .A(n5540), .B(n4409), .Z(n5547) );
  CND2X1 U8047 ( .A(n5534), .B(n4406), .Z(n5541) );
  CND2X1 U8048 ( .A(n5522), .B(n4406), .Z(n5529) );
  CND2X1 U8049 ( .A(n5528), .B(n4408), .Z(n5535) );
  CND2X1 U8050 ( .A(n5466), .B(n4408), .Z(n5470) );
  CND2X1 U8051 ( .A(n5473), .B(n4406), .Z(n5478) );
  CND2X1 U8052 ( .A(n5469), .B(n4406), .Z(n5474) );
  CND2X1 U8053 ( .A(n6555), .B(n4010), .Z(n6565) );
  CANR2X1 U8054 ( .A(N6224), .B(n3594), .C(n3896), .D(n3637), .Z(n2120) );
  CANR2X1 U8055 ( .A(N3109), .B(n3592), .C(N2075), .D(n3637), .Z(n2106) );
  CNIVX1 U8056 ( .A(n79), .Z(n3629) );
  CNIVX1 U8057 ( .A(n79), .Z(n3634) );
  CNIVX1 U8058 ( .A(n79), .Z(n3631) );
  CNIVX1 U8059 ( .A(n79), .Z(n3619) );
  CNIVX1 U8060 ( .A(n79), .Z(n3609) );
  CNIVX1 U8061 ( .A(n79), .Z(n3613) );
  CNIVX1 U8062 ( .A(n79), .Z(n3635) );
  CNIVX1 U8063 ( .A(n79), .Z(n3637) );
  CNIVX1 U8064 ( .A(n79), .Z(n3638) );
  CNIVX1 U8065 ( .A(n73), .Z(n3604) );
  CNIVX1 U8066 ( .A(n73), .Z(n3605) );
  CNIVX1 U8067 ( .A(n4428), .Z(n4001) );
  CNIVX1 U8068 ( .A(n4428), .Z(n3992) );
  CNIVX1 U8069 ( .A(n4428), .Z(n3983) );
  CNIVX1 U8070 ( .A(n4428), .Z(n4002) );
  CNIVX1 U8071 ( .A(n4428), .Z(n3993) );
  CNIVX1 U8072 ( .A(n4428), .Z(n3984) );
  CNIVX1 U8073 ( .A(n4428), .Z(n4004) );
  CNIVX1 U8074 ( .A(n4428), .Z(n3995) );
  CNIVX1 U8075 ( .A(n4428), .Z(n3986) );
  CNIVX1 U8076 ( .A(n4428), .Z(n3996) );
  CNIVX1 U8077 ( .A(n4428), .Z(n3987) );
  CNIVX1 U8078 ( .A(n4428), .Z(n3997) );
  CNIVX1 U8079 ( .A(n4428), .Z(n3988) );
  CNIVX1 U8080 ( .A(n4428), .Z(n3999) );
  CNIVX1 U8081 ( .A(n4428), .Z(n3998) );
  CNIVX1 U8082 ( .A(n4428), .Z(n3990) );
  CNIVX1 U8083 ( .A(n4428), .Z(n3989) );
  CNIVX1 U8084 ( .A(n4428), .Z(n4000) );
  CNIVX1 U8085 ( .A(n4428), .Z(n3991) );
  CNIVX1 U8086 ( .A(n4428), .Z(n3982) );
  CNIVX1 U8087 ( .A(n4428), .Z(n4003) );
  CNIVX1 U8088 ( .A(n4428), .Z(n3994) );
  CNIVX1 U8089 ( .A(n4428), .Z(n3985) );
  CNIVX1 U8090 ( .A(n4428), .Z(n4008) );
  CIVX2 U8091 ( .A(n4295), .Z(n4228) );
  CIVX2 U8092 ( .A(n4295), .Z(n4229) );
  CIVX2 U8093 ( .A(n4295), .Z(n4230) );
  CIVX2 U8094 ( .A(n4295), .Z(n4231) );
  CIVX2 U8095 ( .A(n4295), .Z(n4232) );
  CIVX2 U8096 ( .A(n4295), .Z(n4233) );
  CIVX2 U8097 ( .A(n4295), .Z(n4234) );
  CIVX2 U8098 ( .A(n4295), .Z(n4235) );
  CIVX2 U8099 ( .A(n4295), .Z(n4236) );
  CNIVX1 U8100 ( .A(n4428), .Z(n4007) );
  CNIVX1 U8101 ( .A(n4428), .Z(n4005) );
  CNIVX1 U8102 ( .A(n4428), .Z(n4006) );
  CNIVX1 U8103 ( .A(n4428), .Z(n4009) );
  CND2X1 U8104 ( .A(n6558), .B(n4010), .Z(n6567) );
  CNR2X1 U8105 ( .A(n4439), .B(n15731), .Z(n15734) );
  CNR2X1 U8106 ( .A(n4439), .B(n4440), .Z(n15735) );
  CNR2X1 U8107 ( .A(n4439), .B(n15732), .Z(n15736) );
  CIVX2 U8108 ( .A(n4378), .Z(n4305) );
  CIVX2 U8109 ( .A(n4377), .Z(n4306) );
  CND2X1 U8110 ( .A(n15731), .B(n4439), .Z(n15737) );
  CND2X1 U8111 ( .A(n4439), .B(n4440), .Z(n15738) );
  CND2X1 U8112 ( .A(n4439), .B(n15732), .Z(n15733) );
  CNIVX1 U8113 ( .A(n4415), .Z(n3899) );
  CNIVX1 U8114 ( .A(n4415), .Z(n3928) );
  CNIVX1 U8115 ( .A(n4415), .Z(n3927) );
  CNIVX1 U8116 ( .A(n4415), .Z(n3926) );
  CNIVX1 U8117 ( .A(n4415), .Z(n3925) );
  CNIVX1 U8118 ( .A(n4415), .Z(n3923) );
  CNIVX1 U8119 ( .A(n4415), .Z(n3922) );
  CNIVX1 U8120 ( .A(n4415), .Z(n3921) );
  CNIVX1 U8121 ( .A(n4415), .Z(n3920) );
  CNIVX1 U8122 ( .A(n4415), .Z(n3924) );
  CNIVX1 U8123 ( .A(n4415), .Z(n3939) );
  CNIVX1 U8124 ( .A(n4415), .Z(n3938) );
  CNIVX1 U8125 ( .A(n4415), .Z(n3937) );
  CNIVX1 U8126 ( .A(n4415), .Z(n3936) );
  CNIVX1 U8127 ( .A(n4415), .Z(n3935) );
  CNIVX1 U8128 ( .A(n4415), .Z(n3933) );
  CNIVX1 U8129 ( .A(n4415), .Z(n3932) );
  CNIVX1 U8130 ( .A(n4415), .Z(n3931) );
  CNIVX1 U8131 ( .A(n4415), .Z(n3930) );
  CNIVX1 U8132 ( .A(n4415), .Z(n3929) );
  CNIVX1 U8133 ( .A(n4415), .Z(n3934) );
  CNIVX1 U8134 ( .A(n4415), .Z(n3908) );
  CNIVX1 U8135 ( .A(n4415), .Z(n3907) );
  CNIVX1 U8136 ( .A(n4415), .Z(n3906) );
  CNIVX1 U8137 ( .A(n4415), .Z(n3905) );
  CNIVX1 U8138 ( .A(n4415), .Z(n3903) );
  CNIVX1 U8139 ( .A(n4415), .Z(n3902) );
  CNIVX1 U8140 ( .A(n4415), .Z(n3901) );
  CNIVX1 U8141 ( .A(n4415), .Z(n3900) );
  CNIVX1 U8142 ( .A(n4415), .Z(n3904) );
  CNIVX1 U8143 ( .A(n4415), .Z(n3918) );
  CNIVX1 U8144 ( .A(n4415), .Z(n3917) );
  CNIVX1 U8145 ( .A(n4415), .Z(n3916) );
  CNIVX1 U8146 ( .A(n4415), .Z(n3915) );
  CNIVX1 U8147 ( .A(n4415), .Z(n3913) );
  CNIVX1 U8148 ( .A(n4415), .Z(n3912) );
  CNIVX1 U8149 ( .A(n4415), .Z(n3911) );
  CNIVX1 U8150 ( .A(n4415), .Z(n3910) );
  CNIVX1 U8151 ( .A(n4415), .Z(n3909) );
  CNIVX1 U8152 ( .A(n4415), .Z(n3914) );
  CNIVX1 U8153 ( .A(n4415), .Z(n3919) );
  CNIVX1 U8154 ( .A(n4415), .Z(n3970) );
  CNIVX1 U8155 ( .A(n4415), .Z(n3969) );
  CNIVX1 U8156 ( .A(n4415), .Z(n3968) );
  CNIVX1 U8157 ( .A(n4415), .Z(n3963) );
  CNIVX1 U8158 ( .A(n4415), .Z(n3961) );
  CNIVX1 U8159 ( .A(n4415), .Z(n3979) );
  CNIVX1 U8160 ( .A(n4415), .Z(n3975) );
  CNIVX1 U8161 ( .A(n4415), .Z(n3974) );
  CNIVX1 U8162 ( .A(n4415), .Z(n3973) );
  CNIVX1 U8163 ( .A(n4415), .Z(n3949) );
  CNIVX1 U8164 ( .A(n4415), .Z(n3948) );
  CNIVX1 U8165 ( .A(n4415), .Z(n3947) );
  CNIVX1 U8166 ( .A(n4415), .Z(n3946) );
  CNIVX1 U8167 ( .A(n4415), .Z(n3944) );
  CNIVX1 U8168 ( .A(n4415), .Z(n3943) );
  CNIVX1 U8169 ( .A(n4415), .Z(n3942) );
  CNIVX1 U8170 ( .A(n4415), .Z(n3941) );
  CNIVX1 U8171 ( .A(n4415), .Z(n3940) );
  CNIVX1 U8172 ( .A(n4415), .Z(n3945) );
  CNIVX1 U8173 ( .A(n4415), .Z(n3959) );
  CNIVX1 U8174 ( .A(n4415), .Z(n3958) );
  CNIVX1 U8175 ( .A(n4415), .Z(n3957) );
  CNIVX1 U8176 ( .A(n4415), .Z(n3956) );
  CNIVX1 U8177 ( .A(n4415), .Z(n3954) );
  CNIVX1 U8178 ( .A(n4415), .Z(n3952) );
  CNIVX1 U8179 ( .A(n4415), .Z(n3951) );
  CNIVX1 U8180 ( .A(n4415), .Z(n3960) );
  CNIVX1 U8181 ( .A(n4415), .Z(n3955) );
  CNIVX1 U8182 ( .A(n4415), .Z(n3950) );
  CNIVX1 U8183 ( .A(n4415), .Z(n3967) );
  CNIVX1 U8184 ( .A(n4415), .Z(n3965) );
  CNIVX1 U8185 ( .A(n4415), .Z(n3964) );
  CNIVX1 U8186 ( .A(n4415), .Z(n3966) );
  CNIVX1 U8187 ( .A(n4415), .Z(n3972) );
  CNIVX1 U8188 ( .A(n4415), .Z(n3953) );
  CNIVX1 U8189 ( .A(n4415), .Z(n3980) );
  CNIVX1 U8190 ( .A(n4415), .Z(n3978) );
  CNIVX1 U8191 ( .A(n4415), .Z(n3977) );
  CNIVX1 U8192 ( .A(n4415), .Z(n3971) );
  CNIVX1 U8193 ( .A(n4415), .Z(n3962) );
  CNIVX1 U8194 ( .A(n4415), .Z(n3976) );
  CNIVX1 U8195 ( .A(n4415), .Z(n3981) );
  CEOX1 U8196 ( .A(N766), .B(mem_data1[748]), .Z(N7531) );
  CEOX1 U8197 ( .A(N764), .B(mem_data1[746]), .Z(N7533) );
  CEOX1 U8198 ( .A(N638), .B(mem_data1[620]), .Z(N7659) );
  CEOX1 U8199 ( .A(N636), .B(mem_data1[618]), .Z(N7661) );
  CEOX1 U8200 ( .A(N20), .B(mem_data1[2]), .Z(N8277) );
  CEOX1 U8201 ( .A(N27), .B(mem_data1[9]), .Z(N8270) );
  CNR2X1 U8202 ( .A(n6515), .B(n3834), .Z(N27) );
  CEOX1 U8203 ( .A(N26), .B(mem_data1[8]), .Z(N8271) );
  CNR2X1 U8204 ( .A(n3837), .B(n6398), .Z(N26) );
  CEOX1 U8205 ( .A(N25), .B(mem_data1[7]), .Z(N8272) );
  CEOX1 U8206 ( .A(N24), .B(mem_data1[6]), .Z(N8273) );
  CEOX1 U8207 ( .A(N23), .B(mem_data1[5]), .Z(N8274) );
  CEOX1 U8208 ( .A(N21), .B(mem_data1[3]), .Z(N8276) );
  CEOX1 U8209 ( .A(N19), .B(mem_data1[1]), .Z(N8278) );
  CEOX1 U8210 ( .A(N22), .B(mem_data1[4]), .Z(N8275) );
  CNR2X1 U8211 ( .A(n3853), .B(n5568), .Z(N22) );
  CEOX1 U8212 ( .A(N28), .B(mem_data1[10]), .Z(N8269) );
  CNR2X1 U8213 ( .A(n3835), .B(n4762), .Z(N28) );
  CND2X1 U8214 ( .A(n4816), .B(n3724), .Z(n4567) );
  CEOX1 U8215 ( .A(N31), .B(mem_data1[13]), .Z(N8266) );
  CNR2X1 U8216 ( .A(n3834), .B(n4767), .Z(N31) );
  CEOX1 U8217 ( .A(N30), .B(mem_data1[12]), .Z(N8267) );
  CNR2X1 U8218 ( .A(n3850), .B(n4766), .Z(N30) );
  CEOX1 U8219 ( .A(N29), .B(mem_data1[11]), .Z(N8268) );
  CNR2X1 U8220 ( .A(n3849), .B(n4763), .Z(N29) );
  CND2X1 U8221 ( .A(n4820), .B(n3730), .Z(n4606) );
  CND2X1 U8222 ( .A(n4818), .B(n3724), .Z(n4588) );
  CNR2X1 U8223 ( .A(n3850), .B(n6453), .Z(N112) );
  CEOX1 U8224 ( .A(N18), .B(mem_data1[0]), .Z(N8279) );
  CNR2X1 U8225 ( .A(n3838), .B(n4738), .Z(N18) );
  CEOX1 U8226 ( .A(N466), .B(mem_data1[448]), .Z(N7831) );
  CNR2X1 U8227 ( .A(n3825), .B(n5427), .Z(N466) );
  CEOX1 U8228 ( .A(N1023), .B(mem_data1[1005]), .Z(N7274) );
  CNR2X1 U8229 ( .A(n3817), .B(n6354), .Z(N1023) );
  CEOX1 U8230 ( .A(N1020), .B(mem_data1[1002]), .Z(N7277) );
  CEOX1 U8231 ( .A(N1021), .B(mem_data1[1003]), .Z(N7276) );
  CNR2X1 U8232 ( .A(n3819), .B(n6350), .Z(N1021) );
  CEOX1 U8233 ( .A(N849), .B(mem_data1[831]), .Z(N7448) );
  CEOX1 U8234 ( .A(N772), .B(mem_data1[754]), .Z(N7525) );
  CEOX1 U8235 ( .A(N708), .B(mem_data1[690]), .Z(N7589) );
  CNR2X1 U8236 ( .A(n3823), .B(n5975), .Z(N708) );
  CEOX1 U8237 ( .A(N680), .B(mem_data1[662]), .Z(N7617) );
  CNR2X1 U8238 ( .A(n3829), .B(n5944), .Z(N680) );
  CEOX1 U8239 ( .A(N644), .B(mem_data1[626]), .Z(N7653) );
  CEOX1 U8240 ( .A(N580), .B(mem_data1[562]), .Z(N7717) );
  CNR2X1 U8241 ( .A(n3845), .B(n5975), .Z(N580) );
  CEOX1 U8242 ( .A(N883), .B(mem_data1[865]), .Z(N7414) );
  CEOX1 U8243 ( .A(N552), .B(mem_data1[534]), .Z(N7745) );
  CNR2X1 U8244 ( .A(n3841), .B(n5944), .Z(N552) );
  CEOX1 U8245 ( .A(N1009), .B(mem_data1[991]), .Z(N7288) );
  CNR2X1 U8246 ( .A(n3829), .B(n6503), .Z(N1009) );
  CEOX1 U8247 ( .A(N972), .B(mem_data1[954]), .Z(N7325) );
  CEOX1 U8248 ( .A(N851), .B(mem_data1[833]), .Z(N7446) );
  CNR2X1 U8249 ( .A(n3842), .B(n6466), .Z(N851) );
  CEOX1 U8250 ( .A(N979), .B(mem_data1[961]), .Z(N7318) );
  CNR2X1 U8251 ( .A(n3829), .B(n6466), .Z(N979) );
  CEOX1 U8252 ( .A(N977), .B(mem_data1[959]), .Z(N7320) );
  CEOX1 U8253 ( .A(N915), .B(mem_data1[897]), .Z(N7382) );
  CNR2X1 U8254 ( .A(n3822), .B(n6394), .Z(N915) );
  CEOX1 U8255 ( .A(N787), .B(mem_data1[769]), .Z(N7510) );
  CNR2X1 U8256 ( .A(n3850), .B(n6394), .Z(N787) );
  CEOX1 U8257 ( .A(N793), .B(mem_data1[775]), .Z(N7504) );
  CNR2X1 U8258 ( .A(n3836), .B(n6402), .Z(N793) );
  CEOX1 U8259 ( .A(N751), .B(mem_data1[733]), .Z(N7546) );
  CEOX1 U8260 ( .A(N616), .B(mem_data1[598]), .Z(N7681) );
  CNR2X1 U8261 ( .A(n3852), .B(n6015), .Z(N616) );
  CEOX1 U8262 ( .A(N615), .B(mem_data1[597]), .Z(N7682) );
  CNR2X1 U8263 ( .A(n3851), .B(n6014), .Z(N615) );
  CEOX1 U8264 ( .A(N921), .B(mem_data1[903]), .Z(N7376) );
  CNR2X1 U8265 ( .A(n3821), .B(n6402), .Z(N921) );
  CEOX1 U8266 ( .A(N750), .B(mem_data1[732]), .Z(N7547) );
  CEOX1 U8267 ( .A(N744), .B(mem_data1[726]), .Z(N7553) );
  CNR2X1 U8268 ( .A(n3828), .B(n6015), .Z(N744) );
  CEOX1 U8269 ( .A(N743), .B(mem_data1[725]), .Z(N7554) );
  CNR2X1 U8270 ( .A(n3829), .B(n6014), .Z(N743) );
  CEOX1 U8271 ( .A(N709), .B(mem_data1[691]), .Z(N7588) );
  CNR2X1 U8272 ( .A(n3822), .B(n5976), .Z(N709) );
  CEOX1 U8273 ( .A(N707), .B(mem_data1[689]), .Z(N7590) );
  CNR2X1 U8274 ( .A(n3824), .B(n5973), .Z(N707) );
  CEOX1 U8275 ( .A(N681), .B(mem_data1[663]), .Z(N7616) );
  CNR2X1 U8276 ( .A(n3816), .B(n5945), .Z(N681) );
  CEOX1 U8277 ( .A(N679), .B(mem_data1[661]), .Z(N7618) );
  CNR2X1 U8278 ( .A(n3830), .B(n5943), .Z(N679) );
  CEOX1 U8279 ( .A(N645), .B(mem_data1[627]), .Z(N7652) );
  CEOX1 U8280 ( .A(N643), .B(mem_data1[625]), .Z(N7654) );
  CEOX1 U8281 ( .A(N581), .B(mem_data1[563]), .Z(N7716) );
  CNR2X1 U8282 ( .A(n3846), .B(n5976), .Z(N581) );
  CEOX1 U8283 ( .A(N579), .B(mem_data1[561]), .Z(N7718) );
  CNR2X1 U8284 ( .A(n3844), .B(n5973), .Z(N579) );
  CEOX1 U8285 ( .A(N551), .B(mem_data1[533]), .Z(N7746) );
  CNR2X1 U8286 ( .A(n3840), .B(n5943), .Z(N551) );
  CEOX1 U8287 ( .A(N985), .B(mem_data1[967]), .Z(N7312) );
  CNR2X1 U8288 ( .A(n3828), .B(n6472), .Z(N985) );
  CEOX1 U8289 ( .A(N959), .B(mem_data1[941]), .Z(N7338) );
  CNR2X1 U8290 ( .A(n3826), .B(n6444), .Z(N959) );
  CEOX1 U8291 ( .A(N948), .B(mem_data1[930]), .Z(N7349) );
  CNR2X1 U8292 ( .A(n3833), .B(n6432), .Z(N948) );
  CEOX1 U8293 ( .A(N913), .B(mem_data1[895]), .Z(N7384) );
  CEOX1 U8294 ( .A(N857), .B(mem_data1[839]), .Z(N7440) );
  CNR2X1 U8295 ( .A(n3844), .B(n6472), .Z(N857) );
  CEOX1 U8296 ( .A(N831), .B(mem_data1[813]), .Z(N7466) );
  CNR2X1 U8297 ( .A(n3846), .B(n6444), .Z(N831) );
  CEOX1 U8298 ( .A(N820), .B(mem_data1[802]), .Z(N7477) );
  CNR2X1 U8299 ( .A(n3838), .B(n6432), .Z(N820) );
  CEOX1 U8300 ( .A(N785), .B(mem_data1[767]), .Z(N7512) );
  CEOX1 U8301 ( .A(N971), .B(mem_data1[953]), .Z(N7326) );
  CNR2X1 U8302 ( .A(n3819), .B(n6457), .Z(N971) );
  CEOX1 U8303 ( .A(N947), .B(mem_data1[929]), .Z(N7350) );
  CNR2X1 U8304 ( .A(n3818), .B(n6430), .Z(N947) );
  CEOX1 U8305 ( .A(N819), .B(mem_data1[801]), .Z(N7478) );
  CNR2X1 U8306 ( .A(n3837), .B(n6430), .Z(N819) );
  CEOX1 U8307 ( .A(N522), .B(mem_data1[504]), .Z(N7775) );
  CEOX1 U8308 ( .A(N973), .B(mem_data1[955]), .Z(N7324) );
  CNR2X1 U8309 ( .A(n3815), .B(n6459), .Z(N973) );
  CEOX1 U8310 ( .A(N922), .B(mem_data1[904]), .Z(N7375) );
  CNR2X1 U8311 ( .A(n3826), .B(n6403), .Z(N922) );
  CEOX1 U8312 ( .A(N794), .B(mem_data1[776]), .Z(N7503) );
  CNR2X1 U8313 ( .A(n3837), .B(n6403), .Z(N794) );
  CEOX1 U8314 ( .A(N792), .B(mem_data1[774]), .Z(N7505) );
  CNR2X1 U8315 ( .A(n3835), .B(n6401), .Z(N792) );
  CEOX1 U8316 ( .A(N773), .B(mem_data1[755]), .Z(N7524) );
  CEOX1 U8317 ( .A(N765), .B(mem_data1[747]), .Z(N7532) );
  CEOX1 U8318 ( .A(N749), .B(mem_data1[731]), .Z(N7548) );
  CNR2X1 U8319 ( .A(n3815), .B(n6021), .Z(N749) );
  CEOX1 U8320 ( .A(N701), .B(mem_data1[683]), .Z(N7596) );
  CNR2X1 U8321 ( .A(n3818), .B(n5967), .Z(N701) );
  CEOX1 U8322 ( .A(N637), .B(mem_data1[619]), .Z(N7660) );
  CEOX1 U8323 ( .A(N573), .B(mem_data1[555]), .Z(N7724) );
  CNR2X1 U8324 ( .A(n3842), .B(n5967), .Z(N573) );
  CEOX1 U8325 ( .A(N553), .B(mem_data1[535]), .Z(N7744) );
  CNR2X1 U8326 ( .A(n3842), .B(n5945), .Z(N553) );
  CEOX1 U8327 ( .A(N958), .B(mem_data1[940]), .Z(N7339) );
  CNR2X1 U8328 ( .A(n3825), .B(n6443), .Z(N958) );
  CEOX1 U8329 ( .A(N949), .B(mem_data1[931]), .Z(N7348) );
  CNR2X1 U8330 ( .A(n3825), .B(n6433), .Z(N949) );
  CEOX1 U8331 ( .A(N830), .B(mem_data1[812]), .Z(N7467) );
  CNR2X1 U8332 ( .A(n3845), .B(n6443), .Z(N830) );
  CEOX1 U8333 ( .A(N821), .B(mem_data1[803]), .Z(N7476) );
  CNR2X1 U8334 ( .A(n3851), .B(n6433), .Z(N821) );
  CEOX1 U8335 ( .A(N1008), .B(mem_data1[990]), .Z(N7289) );
  CNR2X1 U8336 ( .A(n3828), .B(n6502), .Z(N1008) );
  CEOX1 U8337 ( .A(N1002), .B(mem_data1[984]), .Z(N7295) );
  CNR2X1 U8338 ( .A(n3827), .B(n6493), .Z(N1002) );
  CEOX1 U8339 ( .A(N1001), .B(mem_data1[983]), .Z(N7296) );
  CEOX1 U8340 ( .A(N984), .B(mem_data1[966]), .Z(N7313) );
  CNR2X1 U8341 ( .A(n3827), .B(n6471), .Z(N984) );
  CEOX1 U8342 ( .A(N920), .B(mem_data1[902]), .Z(N7377) );
  CNR2X1 U8343 ( .A(n3822), .B(n6401), .Z(N920) );
  CEOX1 U8344 ( .A(N884), .B(mem_data1[866]), .Z(N7413) );
  CEOX1 U8345 ( .A(N856), .B(mem_data1[838]), .Z(N7441) );
  CNR2X1 U8346 ( .A(n3843), .B(n6471), .Z(N856) );
  CEOX1 U8347 ( .A(N769), .B(mem_data1[751]), .Z(N7528) );
  CEOX1 U8348 ( .A(N752), .B(mem_data1[734]), .Z(N7545) );
  CNR2X1 U8349 ( .A(n3818), .B(n6024), .Z(N752) );
  CEOX1 U8350 ( .A(N735), .B(mem_data1[717]), .Z(N7562) );
  CNR2X1 U8351 ( .A(n3833), .B(n6005), .Z(N735) );
  CEOX1 U8352 ( .A(N732), .B(mem_data1[714]), .Z(N7565) );
  CNR2X1 U8353 ( .A(n3821), .B(n6002), .Z(N732) );
  CEOX1 U8354 ( .A(N683), .B(mem_data1[665]), .Z(N7614) );
  CNR2X1 U8355 ( .A(n3832), .B(n5947), .Z(N683) );
  CEOX1 U8356 ( .A(N671), .B(mem_data1[653]), .Z(N7626) );
  CNR2X1 U8357 ( .A(n3825), .B(n5934), .Z(N671) );
  CEOX1 U8358 ( .A(N668), .B(mem_data1[650]), .Z(N7629) );
  CNR2X1 U8359 ( .A(n3822), .B(n5931), .Z(N668) );
  CEOX1 U8360 ( .A(N607), .B(mem_data1[589]), .Z(N7690) );
  CNR2X1 U8361 ( .A(n3843), .B(n6005), .Z(N607) );
  CEOX1 U8362 ( .A(N604), .B(mem_data1[586]), .Z(N7693) );
  CNR2X1 U8363 ( .A(n3847), .B(n6002), .Z(N604) );
  CEOX1 U8364 ( .A(N555), .B(mem_data1[537]), .Z(N7742) );
  CNR2X1 U8365 ( .A(n3841), .B(n5947), .Z(N555) );
  CEOX1 U8366 ( .A(N543), .B(mem_data1[525]), .Z(N7754) );
  CNR2X1 U8367 ( .A(n3836), .B(n5934), .Z(N543) );
  CEOX1 U8368 ( .A(N540), .B(mem_data1[522]), .Z(N7757) );
  CNR2X1 U8369 ( .A(n3853), .B(n5931), .Z(N540) );
  CEOX1 U8370 ( .A(N994), .B(mem_data1[976]), .Z(N7303) );
  CNR2X1 U8371 ( .A(n3819), .B(n6482), .Z(N994) );
  CEOX1 U8372 ( .A(N992), .B(mem_data1[974]), .Z(N7305) );
  CNR2X1 U8373 ( .A(n3823), .B(n6480), .Z(N992) );
  CEOX1 U8374 ( .A(N991), .B(mem_data1[973]), .Z(N7306) );
  CNR2X1 U8375 ( .A(n3822), .B(n6479), .Z(N991) );
  CEOX1 U8376 ( .A(N988), .B(mem_data1[970]), .Z(N7309) );
  CNR2X1 U8377 ( .A(n3825), .B(n6476), .Z(N988) );
  CEOX1 U8378 ( .A(N986), .B(mem_data1[968]), .Z(N7311) );
  CNR2X1 U8379 ( .A(n3828), .B(n6473), .Z(N986) );
  CEOX1 U8380 ( .A(N960), .B(mem_data1[942]), .Z(N7337) );
  CNR2X1 U8381 ( .A(n3833), .B(n6445), .Z(N960) );
  CEOX1 U8382 ( .A(N957), .B(mem_data1[939]), .Z(N7340) );
  CNR2X1 U8383 ( .A(n3824), .B(n6441), .Z(N957) );
  CEOX1 U8384 ( .A(N950), .B(mem_data1[932]), .Z(N7347) );
  CNR2X1 U8385 ( .A(n3815), .B(n6434), .Z(N950) );
  CEOX1 U8386 ( .A(N866), .B(mem_data1[848]), .Z(N7431) );
  CNR2X1 U8387 ( .A(n3852), .B(n6482), .Z(N866) );
  CEOX1 U8388 ( .A(N860), .B(mem_data1[842]), .Z(N7437) );
  CNR2X1 U8389 ( .A(n3847), .B(n6476), .Z(N860) );
  CEOX1 U8390 ( .A(N858), .B(mem_data1[840]), .Z(N7439) );
  CNR2X1 U8391 ( .A(n3845), .B(n6473), .Z(N858) );
  CEOX1 U8392 ( .A(N848), .B(mem_data1[830]), .Z(N7449) );
  CNR2X1 U8393 ( .A(n3839), .B(n6462), .Z(N848) );
  CEOX1 U8394 ( .A(N832), .B(mem_data1[814]), .Z(N7465) );
  CNR2X1 U8395 ( .A(n3847), .B(n6445), .Z(N832) );
  CEOX1 U8396 ( .A(N829), .B(mem_data1[811]), .Z(N7468) );
  CNR2X1 U8397 ( .A(n3844), .B(n6441), .Z(N829) );
  CEOX1 U8398 ( .A(N822), .B(mem_data1[804]), .Z(N7475) );
  CNR2X1 U8399 ( .A(n3839), .B(n6434), .Z(N822) );
  CEOX1 U8400 ( .A(N523), .B(mem_data1[505]), .Z(N7774) );
  CEOX1 U8401 ( .A(N521), .B(mem_data1[503]), .Z(N7776) );
  CEOX1 U8402 ( .A(N995), .B(mem_data1[977]), .Z(N7302) );
  CNR2X1 U8403 ( .A(n3820), .B(n6483), .Z(N995) );
  CEOX1 U8404 ( .A(N989), .B(mem_data1[971]), .Z(N7308) );
  CNR2X1 U8405 ( .A(n3826), .B(n6477), .Z(N989) );
  CEOX1 U8406 ( .A(N956), .B(mem_data1[938]), .Z(N7341) );
  CNR2X1 U8407 ( .A(n3829), .B(n6440), .Z(N956) );
  CEOX1 U8408 ( .A(N951), .B(mem_data1[933]), .Z(N7346) );
  CNR2X1 U8409 ( .A(n3830), .B(n6435), .Z(N951) );
  CEOX1 U8410 ( .A(N945), .B(mem_data1[927]), .Z(N7352) );
  CNR2X1 U8411 ( .A(n3816), .B(n6428), .Z(N945) );
  CEOX1 U8412 ( .A(N931), .B(mem_data1[913]), .Z(N7366) );
  CNR2X1 U8413 ( .A(n3833), .B(n6413), .Z(N931) );
  CEOX1 U8414 ( .A(N930), .B(mem_data1[912]), .Z(N7367) );
  CNR2X1 U8415 ( .A(n3830), .B(n6412), .Z(N930) );
  CEOX1 U8416 ( .A(N925), .B(mem_data1[907]), .Z(N7372) );
  CNR2X1 U8417 ( .A(n3829), .B(n6406), .Z(N925) );
  CEOX1 U8418 ( .A(N924), .B(mem_data1[906]), .Z(N7373) );
  CNR2X1 U8419 ( .A(n3824), .B(n6405), .Z(N924) );
  CEOX1 U8420 ( .A(N901), .B(mem_data1[883]), .Z(N7396) );
  CEOX1 U8421 ( .A(N897), .B(mem_data1[879]), .Z(N7400) );
  CEOX1 U8422 ( .A(N881), .B(mem_data1[863]), .Z(N7416) );
  CNR2X1 U8423 ( .A(n3851), .B(n6503), .Z(N881) );
  CEOX1 U8424 ( .A(N867), .B(mem_data1[849]), .Z(N7430) );
  CNR2X1 U8425 ( .A(n3853), .B(n6483), .Z(N867) );
  CEOX1 U8426 ( .A(N861), .B(mem_data1[843]), .Z(N7436) );
  CNR2X1 U8427 ( .A(n3848), .B(n6477), .Z(N861) );
  CEOX1 U8428 ( .A(N852), .B(mem_data1[834]), .Z(N7445) );
  CNR2X1 U8429 ( .A(n3843), .B(n6467), .Z(N852) );
  CEOX1 U8430 ( .A(N828), .B(mem_data1[810]), .Z(N7469) );
  CNR2X1 U8431 ( .A(n3843), .B(n6440), .Z(N828) );
  CEOX1 U8432 ( .A(N823), .B(mem_data1[805]), .Z(N7474) );
  CNR2X1 U8433 ( .A(n3838), .B(n6435), .Z(N823) );
  CEOX1 U8434 ( .A(N817), .B(mem_data1[799]), .Z(N7480) );
  CNR2X1 U8435 ( .A(n3836), .B(n6428), .Z(N817) );
  CEOX1 U8436 ( .A(N803), .B(mem_data1[785]), .Z(N7494) );
  CNR2X1 U8437 ( .A(n3850), .B(n6413), .Z(N803) );
  CEOX1 U8438 ( .A(N802), .B(mem_data1[784]), .Z(N7495) );
  CNR2X1 U8439 ( .A(n3835), .B(n6412), .Z(N802) );
  CEOX1 U8440 ( .A(N800), .B(mem_data1[782]), .Z(N7497) );
  CNR2X1 U8441 ( .A(n3850), .B(n6410), .Z(N800) );
  CEOX1 U8442 ( .A(N799), .B(mem_data1[781]), .Z(N7498) );
  CNR2X1 U8443 ( .A(n3843), .B(n6408), .Z(N799) );
  CEOX1 U8444 ( .A(N797), .B(mem_data1[779]), .Z(N7500) );
  CNR2X1 U8445 ( .A(n3840), .B(n6406), .Z(N797) );
  CEOX1 U8446 ( .A(N796), .B(mem_data1[778]), .Z(N7501) );
  CNR2X1 U8447 ( .A(n3839), .B(n6405), .Z(N796) );
  CEOX1 U8448 ( .A(N767), .B(mem_data1[749]), .Z(N7530) );
  CEOX1 U8449 ( .A(N763), .B(mem_data1[745]), .Z(N7534) );
  CEOX1 U8450 ( .A(N761), .B(mem_data1[743]), .Z(N7536) );
  CEOX1 U8451 ( .A(N759), .B(mem_data1[741]), .Z(N7538) );
  CEOX1 U8452 ( .A(N755), .B(mem_data1[737]), .Z(N7542) );
  CEOX1 U8453 ( .A(N753), .B(mem_data1[735]), .Z(N7544) );
  CNR2X1 U8454 ( .A(n3817), .B(n6025), .Z(N753) );
  CEOX1 U8455 ( .A(N747), .B(mem_data1[729]), .Z(N7550) );
  CNR2X1 U8456 ( .A(n3831), .B(n6018), .Z(N747) );
  CEOX1 U8457 ( .A(N745), .B(mem_data1[727]), .Z(N7552) );
  CNR2X1 U8458 ( .A(n3833), .B(n6016), .Z(N745) );
  CEOX1 U8459 ( .A(N742), .B(mem_data1[724]), .Z(N7555) );
  CNR2X1 U8460 ( .A(n3830), .B(n6013), .Z(N742) );
  CEOX1 U8461 ( .A(N739), .B(mem_data1[721]), .Z(N7558) );
  CNR2X1 U8462 ( .A(n3827), .B(n6010), .Z(N739) );
  CEOX1 U8463 ( .A(N737), .B(mem_data1[719]), .Z(N7560) );
  CNR2X1 U8464 ( .A(n3829), .B(n6007), .Z(N737) );
  CEOX1 U8465 ( .A(N703), .B(mem_data1[685]), .Z(N7594) );
  CNR2X1 U8466 ( .A(n3816), .B(n5969), .Z(N703) );
  CEOX1 U8467 ( .A(N699), .B(mem_data1[681]), .Z(N7598) );
  CNR2X1 U8468 ( .A(n3826), .B(n5965), .Z(N699) );
  CEOX1 U8469 ( .A(N697), .B(mem_data1[679]), .Z(N7600) );
  CNR2X1 U8470 ( .A(n3819), .B(n5962), .Z(N697) );
  CEOX1 U8471 ( .A(N695), .B(mem_data1[677]), .Z(N7602) );
  CNR2X1 U8472 ( .A(n3823), .B(n5960), .Z(N695) );
  CEOX1 U8473 ( .A(N691), .B(mem_data1[673]), .Z(N7606) );
  CNR2X1 U8474 ( .A(n3829), .B(n5956), .Z(N691) );
  CEOX1 U8475 ( .A(N689), .B(mem_data1[671]), .Z(N7608) );
  CNR2X1 U8476 ( .A(n3831), .B(n5954), .Z(N689) );
  CEOX1 U8477 ( .A(N675), .B(mem_data1[657]), .Z(N7622) );
  CNR2X1 U8478 ( .A(n3827), .B(n5938), .Z(N675) );
  CEOX1 U8479 ( .A(N673), .B(mem_data1[655]), .Z(N7624) );
  CNR2X1 U8480 ( .A(n3820), .B(n5936), .Z(N673) );
  CEOX1 U8481 ( .A(N663), .B(mem_data1[645]), .Z(N7634) );
  CNR2X1 U8482 ( .A(n3815), .B(n5925), .Z(N663) );
  CEOX1 U8483 ( .A(N661), .B(mem_data1[643]), .Z(N7636) );
  CNR2X1 U8484 ( .A(n3817), .B(n5923), .Z(N661) );
  CEOX1 U8485 ( .A(N639), .B(mem_data1[621]), .Z(N7658) );
  CEOX1 U8486 ( .A(N635), .B(mem_data1[617]), .Z(N7662) );
  CEOX1 U8487 ( .A(N633), .B(mem_data1[615]), .Z(N7664) );
  CEOX1 U8488 ( .A(N631), .B(mem_data1[613]), .Z(N7666) );
  CEOX1 U8489 ( .A(N627), .B(mem_data1[609]), .Z(N7670) );
  CEOX1 U8490 ( .A(N625), .B(mem_data1[607]), .Z(N7672) );
  CNR2X1 U8491 ( .A(n3837), .B(n6025), .Z(N625) );
  CEOX1 U8492 ( .A(N624), .B(mem_data1[606]), .Z(N7673) );
  CNR2X1 U8493 ( .A(n3836), .B(n6024), .Z(N624) );
  CEOX1 U8494 ( .A(N622), .B(mem_data1[604]), .Z(N7675) );
  CNR2X1 U8495 ( .A(n3848), .B(n6022), .Z(N622) );
  CEOX1 U8496 ( .A(N621), .B(mem_data1[603]), .Z(N7676) );
  CNR2X1 U8497 ( .A(n3849), .B(n6021), .Z(N621) );
  CEOX1 U8498 ( .A(N619), .B(mem_data1[601]), .Z(N7678) );
  CNR2X1 U8499 ( .A(n3848), .B(n6018), .Z(N619) );
  CEOX1 U8500 ( .A(N617), .B(mem_data1[599]), .Z(N7680) );
  CNR2X1 U8501 ( .A(n3853), .B(n6016), .Z(N617) );
  CEOX1 U8502 ( .A(N614), .B(mem_data1[596]), .Z(N7683) );
  CNR2X1 U8503 ( .A(n3850), .B(n6013), .Z(N614) );
  CEOX1 U8504 ( .A(N611), .B(mem_data1[593]), .Z(N7686) );
  CNR2X1 U8505 ( .A(n3847), .B(n6010), .Z(N611) );
  CEOX1 U8506 ( .A(N609), .B(mem_data1[591]), .Z(N7688) );
  CNR2X1 U8507 ( .A(n3844), .B(n6007), .Z(N609) );
  CEOX1 U8508 ( .A(N595), .B(mem_data1[577]), .Z(N7702) );
  CNR2X1 U8509 ( .A(n3835), .B(n5992), .Z(N595) );
  CEOX1 U8510 ( .A(N593), .B(mem_data1[575]), .Z(N7704) );
  CNR2X1 U8511 ( .A(n3853), .B(n5990), .Z(N593) );
  CEOX1 U8512 ( .A(N575), .B(mem_data1[557]), .Z(N7722) );
  CNR2X1 U8513 ( .A(n3839), .B(n5969), .Z(N575) );
  CEOX1 U8514 ( .A(N571), .B(mem_data1[553]), .Z(N7726) );
  CNR2X1 U8515 ( .A(n3836), .B(n5965), .Z(N571) );
  CEOX1 U8516 ( .A(N569), .B(mem_data1[551]), .Z(N7728) );
  CNR2X1 U8517 ( .A(n3834), .B(n5962), .Z(N569) );
  CEOX1 U8518 ( .A(N567), .B(mem_data1[549]), .Z(N7730) );
  CNR2X1 U8519 ( .A(n3840), .B(n5960), .Z(N567) );
  CEOX1 U8520 ( .A(N563), .B(mem_data1[545]), .Z(N7734) );
  CNR2X1 U8521 ( .A(n3852), .B(n5956), .Z(N563) );
  CEOX1 U8522 ( .A(N561), .B(mem_data1[543]), .Z(N7736) );
  CNR2X1 U8523 ( .A(n3850), .B(n5954), .Z(N561) );
  CEOX1 U8524 ( .A(N547), .B(mem_data1[529]), .Z(N7750) );
  CNR2X1 U8525 ( .A(n3844), .B(n5938), .Z(N547) );
  CEOX1 U8526 ( .A(N545), .B(mem_data1[527]), .Z(N7752) );
  CNR2X1 U8527 ( .A(n3838), .B(n5936), .Z(N545) );
  CEOX1 U8528 ( .A(N535), .B(mem_data1[517]), .Z(N7762) );
  CNR2X1 U8529 ( .A(n3848), .B(n5925), .Z(N535) );
  CEOX1 U8530 ( .A(N533), .B(mem_data1[515]), .Z(N7764) );
  CNR2X1 U8531 ( .A(n3846), .B(n5923), .Z(N533) );
  CEOX1 U8532 ( .A(N531), .B(mem_data1[513]), .Z(N7766) );
  CNR2X1 U8533 ( .A(n3843), .B(n5921), .Z(N531) );
  CEOX1 U8534 ( .A(N529), .B(mem_data1[511]), .Z(N7768) );
  CEOX1 U8535 ( .A(N980), .B(mem_data1[962]), .Z(N7317) );
  CNR2X1 U8536 ( .A(n3830), .B(n6467), .Z(N980) );
  CEOX1 U8537 ( .A(N976), .B(mem_data1[958]), .Z(N7321) );
  CNR2X1 U8538 ( .A(n3832), .B(n6462), .Z(N976) );
  CEOX1 U8539 ( .A(N916), .B(mem_data1[898]), .Z(N7381) );
  CNR2X1 U8540 ( .A(n3820), .B(n6395), .Z(N916) );
  CEOX1 U8541 ( .A(N864), .B(mem_data1[846]), .Z(N7433) );
  CNR2X1 U8542 ( .A(n3850), .B(n6480), .Z(N864) );
  CEOX1 U8543 ( .A(N863), .B(mem_data1[845]), .Z(N7434) );
  CNR2X1 U8544 ( .A(n3850), .B(n6479), .Z(N863) );
  CEOX1 U8545 ( .A(N788), .B(mem_data1[770]), .Z(N7509) );
  CNR2X1 U8546 ( .A(n3852), .B(n6395), .Z(N788) );
  CEOX1 U8547 ( .A(N1007), .B(mem_data1[989]), .Z(N7290) );
  CNR2X1 U8548 ( .A(n3833), .B(n6498), .Z(N1007) );
  CEOX1 U8549 ( .A(N928), .B(mem_data1[910]), .Z(N7369) );
  CNR2X1 U8550 ( .A(n3832), .B(n6410), .Z(N928) );
  CEOX1 U8551 ( .A(N927), .B(mem_data1[909]), .Z(N7370) );
  CNR2X1 U8552 ( .A(n3827), .B(n6408), .Z(N927) );
  CEOX1 U8553 ( .A(N902), .B(mem_data1[884]), .Z(N7395) );
  CEOX1 U8554 ( .A(N900), .B(mem_data1[882]), .Z(N7397) );
  CEOX1 U8555 ( .A(N898), .B(mem_data1[880]), .Z(N7399) );
  CEOX1 U8556 ( .A(N896), .B(mem_data1[878]), .Z(N7401) );
  CEOX1 U8557 ( .A(N885), .B(mem_data1[867]), .Z(N7412) );
  CEOX1 U8558 ( .A(N774), .B(mem_data1[756]), .Z(N7523) );
  CEOX1 U8559 ( .A(N768), .B(mem_data1[750]), .Z(N7529) );
  CEOX1 U8560 ( .A(N736), .B(mem_data1[718]), .Z(N7561) );
  CNR2X1 U8561 ( .A(n3824), .B(n6006), .Z(N736) );
  CEOX1 U8562 ( .A(N731), .B(mem_data1[713]), .Z(N7566) );
  CNR2X1 U8563 ( .A(n3822), .B(n6001), .Z(N731) );
  CEOX1 U8564 ( .A(N687), .B(mem_data1[669]), .Z(N7610) );
  CNR2X1 U8565 ( .A(n3827), .B(n5951), .Z(N687) );
  CEOX1 U8566 ( .A(N686), .B(mem_data1[668]), .Z(N7611) );
  CNR2X1 U8567 ( .A(n3818), .B(n5950), .Z(N686) );
  CEOX1 U8568 ( .A(N682), .B(mem_data1[664]), .Z(N7615) );
  CNR2X1 U8569 ( .A(n3833), .B(n5946), .Z(N682) );
  CEOX1 U8570 ( .A(N672), .B(mem_data1[654]), .Z(N7625) );
  CNR2X1 U8571 ( .A(n3824), .B(n5935), .Z(N672) );
  CEOX1 U8572 ( .A(N667), .B(mem_data1[649]), .Z(N7630) );
  CNR2X1 U8573 ( .A(n3823), .B(n5929), .Z(N667) );
  CEOX1 U8574 ( .A(N608), .B(mem_data1[590]), .Z(N7689) );
  CNR2X1 U8575 ( .A(n3845), .B(n6006), .Z(N608) );
  CEOX1 U8576 ( .A(N603), .B(mem_data1[585]), .Z(N7694) );
  CNR2X1 U8577 ( .A(n3846), .B(n6001), .Z(N603) );
  CEOX1 U8578 ( .A(N559), .B(mem_data1[541]), .Z(N7738) );
  CNR2X1 U8579 ( .A(n3848), .B(n5951), .Z(N559) );
  CEOX1 U8580 ( .A(N558), .B(mem_data1[540]), .Z(N7739) );
  CNR2X1 U8581 ( .A(n3847), .B(n5950), .Z(N558) );
  CEOX1 U8582 ( .A(N554), .B(mem_data1[536]), .Z(N7743) );
  CNR2X1 U8583 ( .A(n3843), .B(n5946), .Z(N554) );
  CEOX1 U8584 ( .A(N544), .B(mem_data1[526]), .Z(N7753) );
  CNR2X1 U8585 ( .A(n3837), .B(n5935), .Z(N544) );
  CEOX1 U8586 ( .A(N539), .B(mem_data1[521]), .Z(N7758) );
  CNR2X1 U8587 ( .A(n3852), .B(n5929), .Z(N539) );
  CEOX1 U8588 ( .A(N1006), .B(mem_data1[988]), .Z(N7291) );
  CNR2X1 U8589 ( .A(n3832), .B(n6497), .Z(N1006) );
  CEOX1 U8590 ( .A(N993), .B(mem_data1[975]), .Z(N7304) );
  CNR2X1 U8591 ( .A(n3818), .B(n6481), .Z(N993) );
  CEOX1 U8592 ( .A(N987), .B(mem_data1[969]), .Z(N7310) );
  CNR2X1 U8593 ( .A(n3824), .B(n6474), .Z(N987) );
  CEOX1 U8594 ( .A(N912), .B(mem_data1[894]), .Z(N7385) );
  CEOX1 U8595 ( .A(N886), .B(mem_data1[868]), .Z(N7411) );
  CEOX1 U8596 ( .A(N865), .B(mem_data1[847]), .Z(N7432) );
  CNR2X1 U8597 ( .A(n3851), .B(n6481), .Z(N865) );
  CEOX1 U8598 ( .A(N859), .B(mem_data1[841]), .Z(N7438) );
  CNR2X1 U8599 ( .A(n3846), .B(n6474), .Z(N859) );
  CEOX1 U8600 ( .A(N784), .B(mem_data1[766]), .Z(N7513) );
  CEOX1 U8601 ( .A(N775), .B(mem_data1[757]), .Z(N7522) );
  CEOX1 U8602 ( .A(N520), .B(mem_data1[502]), .Z(N7777) );
  CEOX1 U8603 ( .A(N365), .B(mem_data1[347]), .Z(N7932) );
  CNR2X1 U8604 ( .A(n3851), .B(n5457), .Z(N365) );
  CEOX1 U8605 ( .A(N1005), .B(mem_data1[987]), .Z(N7292) );
  CNR2X1 U8606 ( .A(n3831), .B(n6496), .Z(N1005) );
  CEOX1 U8607 ( .A(N1004), .B(mem_data1[986]), .Z(N7293) );
  CNR2X1 U8608 ( .A(n3831), .B(n6495), .Z(N1004) );
  CEOX1 U8609 ( .A(N1003), .B(mem_data1[985]), .Z(N7294) );
  CNR2X1 U8610 ( .A(n3815), .B(n6494), .Z(N1003) );
  CEOX1 U8611 ( .A(N1000), .B(mem_data1[982]), .Z(N7297) );
  CNR2X1 U8612 ( .A(n3823), .B(n6491), .Z(N1000) );
  CEOX1 U8613 ( .A(N999), .B(mem_data1[981]), .Z(N7298) );
  CNR2X1 U8614 ( .A(n3819), .B(n6490), .Z(N999) );
  CEOX1 U8615 ( .A(N998), .B(mem_data1[980]), .Z(N7299) );
  CNR2X1 U8616 ( .A(n3817), .B(n6489), .Z(N998) );
  CEOX1 U8617 ( .A(N997), .B(mem_data1[979]), .Z(N7300) );
  CNR2X1 U8618 ( .A(n3816), .B(n6485), .Z(N997) );
  CEOX1 U8619 ( .A(N996), .B(mem_data1[978]), .Z(N7301) );
  CNR2X1 U8620 ( .A(n3815), .B(n6484), .Z(N996) );
  CEOX1 U8621 ( .A(N990), .B(mem_data1[972]), .Z(N7307) );
  CNR2X1 U8622 ( .A(n3821), .B(n6478), .Z(N990) );
  CEOX1 U8623 ( .A(N983), .B(mem_data1[965]), .Z(N7314) );
  CNR2X1 U8624 ( .A(n3820), .B(n6470), .Z(N983) );
  CEOX1 U8625 ( .A(N982), .B(mem_data1[964]), .Z(N7315) );
  CNR2X1 U8626 ( .A(n3832), .B(n6469), .Z(N982) );
  CEOX1 U8627 ( .A(N981), .B(mem_data1[963]), .Z(N7316) );
  CNR2X1 U8628 ( .A(n3816), .B(n6468), .Z(N981) );
  CEOX1 U8629 ( .A(N975), .B(mem_data1[957]), .Z(N7322) );
  CNR2X1 U8630 ( .A(n3831), .B(n6461), .Z(N975) );
  CEOX1 U8631 ( .A(N974), .B(mem_data1[956]), .Z(N7323) );
  CNR2X1 U8632 ( .A(n3816), .B(n6460), .Z(N974) );
  CEOX1 U8633 ( .A(N970), .B(mem_data1[952]), .Z(N7327) );
  CNR2X1 U8634 ( .A(n3818), .B(n6456), .Z(N970) );
  CEOX1 U8635 ( .A(N969), .B(mem_data1[951]), .Z(N7328) );
  CNR2X1 U8636 ( .A(n3817), .B(n6455), .Z(N969) );
  CEOX1 U8637 ( .A(N968), .B(mem_data1[950]), .Z(N7329) );
  CNR2X1 U8638 ( .A(n3822), .B(n6454), .Z(N968) );
  CEOX1 U8639 ( .A(N967), .B(mem_data1[949]), .Z(N7330) );
  CNR2X1 U8640 ( .A(n3821), .B(n6452), .Z(N967) );
  CEOX1 U8641 ( .A(N966), .B(mem_data1[948]), .Z(N7331) );
  CNR2X1 U8642 ( .A(n3820), .B(n6451), .Z(N966) );
  CEOX1 U8643 ( .A(N965), .B(mem_data1[947]), .Z(N7332) );
  CNR2X1 U8644 ( .A(n3817), .B(n6450), .Z(N965) );
  CEOX1 U8645 ( .A(N964), .B(mem_data1[946]), .Z(N7333) );
  CNR2X1 U8646 ( .A(n3829), .B(n6449), .Z(N964) );
  CEOX1 U8647 ( .A(N963), .B(mem_data1[945]), .Z(N7334) );
  CNR2X1 U8648 ( .A(n3823), .B(n6448), .Z(N963) );
  CEOX1 U8649 ( .A(N962), .B(mem_data1[944]), .Z(N7335) );
  CNR2X1 U8650 ( .A(n3825), .B(n6447), .Z(N962) );
  CEOX1 U8651 ( .A(N961), .B(mem_data1[943]), .Z(N7336) );
  CNR2X1 U8652 ( .A(n3821), .B(n6446), .Z(N961) );
  CEOX1 U8653 ( .A(N955), .B(mem_data1[937]), .Z(N7342) );
  CNR2X1 U8654 ( .A(n3828), .B(n6439), .Z(N955) );
  CEOX1 U8655 ( .A(N954), .B(mem_data1[936]), .Z(N7343) );
  CNR2X1 U8656 ( .A(n3827), .B(n6438), .Z(N954) );
  CEOX1 U8657 ( .A(N953), .B(mem_data1[935]), .Z(N7344) );
  CNR2X1 U8658 ( .A(n3832), .B(n6437), .Z(N953) );
  CEOX1 U8659 ( .A(N952), .B(mem_data1[934]), .Z(N7345) );
  CNR2X1 U8660 ( .A(n3831), .B(n6436), .Z(N952) );
  CEOX1 U8661 ( .A(N944), .B(mem_data1[926]), .Z(N7353) );
  CNR2X1 U8662 ( .A(n3830), .B(n6427), .Z(N944) );
  CEOX1 U8663 ( .A(N943), .B(mem_data1[925]), .Z(N7354) );
  CNR2X1 U8664 ( .A(n3818), .B(n6426), .Z(N943) );
  CEOX1 U8665 ( .A(N942), .B(mem_data1[924]), .Z(N7355) );
  CNR2X1 U8666 ( .A(n3830), .B(n6425), .Z(N942) );
  CEOX1 U8667 ( .A(N941), .B(mem_data1[923]), .Z(N7356) );
  CNR2X1 U8668 ( .A(n3819), .B(n6424), .Z(N941) );
  CEOX1 U8669 ( .A(N940), .B(mem_data1[922]), .Z(N7357) );
  CNR2X1 U8670 ( .A(n3826), .B(n6423), .Z(N940) );
  CEOX1 U8671 ( .A(N939), .B(mem_data1[921]), .Z(N7358) );
  CNR2X1 U8672 ( .A(n3822), .B(n6422), .Z(N939) );
  CEOX1 U8673 ( .A(N938), .B(mem_data1[920]), .Z(N7359) );
  CNR2X1 U8674 ( .A(n3822), .B(n6421), .Z(N938) );
  CEOX1 U8675 ( .A(N937), .B(mem_data1[919]), .Z(N7360) );
  CNR2X1 U8676 ( .A(n3821), .B(n6419), .Z(N937) );
  CEOX1 U8677 ( .A(N936), .B(mem_data1[918]), .Z(N7361) );
  CNR2X1 U8678 ( .A(n3820), .B(n6418), .Z(N936) );
  CEOX1 U8679 ( .A(N935), .B(mem_data1[917]), .Z(N7362) );
  CNR2X1 U8680 ( .A(n3825), .B(n6417), .Z(N935) );
  CEOX1 U8681 ( .A(N934), .B(mem_data1[916]), .Z(N7363) );
  CNR2X1 U8682 ( .A(n3824), .B(n6416), .Z(N934) );
  CEOX1 U8683 ( .A(N933), .B(mem_data1[915]), .Z(N7364) );
  CNR2X1 U8684 ( .A(n3823), .B(n6415), .Z(N933) );
  CEOX1 U8685 ( .A(N932), .B(mem_data1[914]), .Z(N7365) );
  CNR2X1 U8686 ( .A(n3828), .B(n6414), .Z(N932) );
  CEOX1 U8687 ( .A(N929), .B(mem_data1[911]), .Z(N7368) );
  CNR2X1 U8688 ( .A(n3831), .B(n6411), .Z(N929) );
  CEOX1 U8689 ( .A(N926), .B(mem_data1[908]), .Z(N7371) );
  CNR2X1 U8690 ( .A(n3828), .B(n6407), .Z(N926) );
  CEOX1 U8691 ( .A(N923), .B(mem_data1[905]), .Z(N7374) );
  CNR2X1 U8692 ( .A(n3825), .B(n6404), .Z(N923) );
  CEOX1 U8693 ( .A(N919), .B(mem_data1[901]), .Z(N7378) );
  CNR2X1 U8694 ( .A(n3823), .B(n6400), .Z(N919) );
  CEOX1 U8695 ( .A(N918), .B(mem_data1[900]), .Z(N7379) );
  CNR2X1 U8696 ( .A(n3830), .B(n6399), .Z(N918) );
  CEOX1 U8697 ( .A(N917), .B(mem_data1[899]), .Z(N7380) );
  CNR2X1 U8698 ( .A(n3819), .B(n6396), .Z(N917) );
  CEOX1 U8699 ( .A(N911), .B(mem_data1[893]), .Z(N7386) );
  CEOX1 U8700 ( .A(N910), .B(mem_data1[892]), .Z(N7387) );
  CEOX1 U8701 ( .A(N909), .B(mem_data1[891]), .Z(N7388) );
  CEOX1 U8702 ( .A(N908), .B(mem_data1[890]), .Z(N7389) );
  CEOX1 U8703 ( .A(N907), .B(mem_data1[889]), .Z(N7390) );
  CEOX1 U8704 ( .A(N906), .B(mem_data1[888]), .Z(N7391) );
  CEOX1 U8705 ( .A(N905), .B(mem_data1[887]), .Z(N7392) );
  CEOX1 U8706 ( .A(N904), .B(mem_data1[886]), .Z(N7393) );
  CEOX1 U8707 ( .A(N903), .B(mem_data1[885]), .Z(N7394) );
  CEOX1 U8708 ( .A(N899), .B(mem_data1[881]), .Z(N7398) );
  CEOX1 U8709 ( .A(N895), .B(mem_data1[877]), .Z(N7402) );
  CEOX1 U8710 ( .A(N894), .B(mem_data1[876]), .Z(N7403) );
  CEOX1 U8711 ( .A(N893), .B(mem_data1[875]), .Z(N7404) );
  CEOX1 U8712 ( .A(N892), .B(mem_data1[874]), .Z(N7405) );
  CEOX1 U8713 ( .A(N891), .B(mem_data1[873]), .Z(N7406) );
  CEOX1 U8714 ( .A(N890), .B(mem_data1[872]), .Z(N7407) );
  CEOX1 U8715 ( .A(N889), .B(mem_data1[871]), .Z(N7408) );
  CEOX1 U8716 ( .A(N888), .B(mem_data1[870]), .Z(N7409) );
  CEOX1 U8717 ( .A(N887), .B(mem_data1[869]), .Z(N7410) );
  CEOX1 U8718 ( .A(N880), .B(mem_data1[862]), .Z(N7417) );
  CNR2X1 U8719 ( .A(n3843), .B(n6502), .Z(N880) );
  CEOX1 U8720 ( .A(N879), .B(mem_data1[861]), .Z(N7418) );
  CNR2X1 U8721 ( .A(n3842), .B(n6498), .Z(N879) );
  CEOX1 U8722 ( .A(N878), .B(mem_data1[860]), .Z(N7419) );
  CNR2X1 U8723 ( .A(n3841), .B(n6497), .Z(N878) );
  CEOX1 U8724 ( .A(N877), .B(mem_data1[859]), .Z(N7420) );
  CNR2X1 U8725 ( .A(n3848), .B(n6496), .Z(N877) );
  CEOX1 U8726 ( .A(N876), .B(mem_data1[858]), .Z(N7421) );
  CNR2X1 U8727 ( .A(n3834), .B(n6495), .Z(N876) );
  CEOX1 U8728 ( .A(N875), .B(mem_data1[857]), .Z(N7422) );
  CNR2X1 U8729 ( .A(n3847), .B(n6494), .Z(N875) );
  CEOX1 U8730 ( .A(N874), .B(mem_data1[856]), .Z(N7423) );
  CNR2X1 U8731 ( .A(n3846), .B(n6493), .Z(N874) );
  CEOX1 U8732 ( .A(N873), .B(mem_data1[855]), .Z(N7424) );
  CNR2X1 U8733 ( .A(n3834), .B(n6492), .Z(N873) );
  CEOX1 U8734 ( .A(N872), .B(mem_data1[854]), .Z(N7425) );
  CNR2X1 U8735 ( .A(n3839), .B(n6491), .Z(N872) );
  CEOX1 U8736 ( .A(N871), .B(mem_data1[853]), .Z(N7426) );
  CNR2X1 U8737 ( .A(n3838), .B(n6490), .Z(N871) );
  CEOX1 U8738 ( .A(N870), .B(mem_data1[852]), .Z(N7427) );
  CNR2X1 U8739 ( .A(n3837), .B(n6489), .Z(N870) );
  CEOX1 U8740 ( .A(N869), .B(mem_data1[851]), .Z(N7428) );
  CNR2X1 U8741 ( .A(n3836), .B(n6485), .Z(N869) );
  CEOX1 U8742 ( .A(N868), .B(mem_data1[850]), .Z(N7429) );
  CNR2X1 U8743 ( .A(n3835), .B(n6484), .Z(N868) );
  CEOX1 U8744 ( .A(N862), .B(mem_data1[844]), .Z(N7435) );
  CNR2X1 U8745 ( .A(n3849), .B(n6478), .Z(N862) );
  CEOX1 U8746 ( .A(N855), .B(mem_data1[837]), .Z(N7442) );
  CNR2X1 U8747 ( .A(n3853), .B(n6470), .Z(N855) );
  CEOX1 U8748 ( .A(N854), .B(mem_data1[836]), .Z(N7443) );
  CNR2X1 U8749 ( .A(n3845), .B(n6469), .Z(N854) );
  CEOX1 U8750 ( .A(N853), .B(mem_data1[835]), .Z(N7444) );
  CNR2X1 U8751 ( .A(n3844), .B(n6468), .Z(N853) );
  CEOX1 U8752 ( .A(N847), .B(mem_data1[829]), .Z(N7450) );
  CNR2X1 U8753 ( .A(n3837), .B(n6461), .Z(N847) );
  CEOX1 U8754 ( .A(N846), .B(mem_data1[828]), .Z(N7451) );
  CNR2X1 U8755 ( .A(n3836), .B(n6460), .Z(N846) );
  CEOX1 U8756 ( .A(N845), .B(mem_data1[827]), .Z(N7452) );
  CNR2X1 U8757 ( .A(n3849), .B(n6459), .Z(N845) );
  CEOX1 U8758 ( .A(N844), .B(mem_data1[826]), .Z(N7453) );
  CNR2X1 U8759 ( .A(n3835), .B(n6458), .Z(N844) );
  CEOX1 U8760 ( .A(N843), .B(mem_data1[825]), .Z(N7454) );
  CNR2X1 U8761 ( .A(n3834), .B(n6457), .Z(N843) );
  CEOX1 U8762 ( .A(N842), .B(mem_data1[824]), .Z(N7455) );
  CNR2X1 U8763 ( .A(n3853), .B(n6456), .Z(N842) );
  CEOX1 U8764 ( .A(N841), .B(mem_data1[823]), .Z(N7456) );
  CNR2X1 U8765 ( .A(n3852), .B(n6455), .Z(N841) );
  CEOX1 U8766 ( .A(N840), .B(mem_data1[822]), .Z(N7457) );
  CNR2X1 U8767 ( .A(n3842), .B(n6454), .Z(N840) );
  CEOX1 U8768 ( .A(N839), .B(mem_data1[821]), .Z(N7458) );
  CNR2X1 U8769 ( .A(n3852), .B(n6452), .Z(N839) );
  CEOX1 U8770 ( .A(N838), .B(mem_data1[820]), .Z(N7459) );
  CNR2X1 U8771 ( .A(n3841), .B(n6451), .Z(N838) );
  CEOX1 U8772 ( .A(N837), .B(mem_data1[819]), .Z(N7460) );
  CNR2X1 U8773 ( .A(n3852), .B(n6450), .Z(N837) );
  CEOX1 U8774 ( .A(N836), .B(mem_data1[818]), .Z(N7461) );
  CNR2X1 U8775 ( .A(n3851), .B(n6449), .Z(N836) );
  CEOX1 U8776 ( .A(N835), .B(mem_data1[817]), .Z(N7462) );
  CNR2X1 U8777 ( .A(n3850), .B(n6448), .Z(N835) );
  CEOX1 U8778 ( .A(N834), .B(mem_data1[816]), .Z(N7463) );
  CNR2X1 U8779 ( .A(n3849), .B(n6447), .Z(N834) );
  CEOX1 U8780 ( .A(N833), .B(mem_data1[815]), .Z(N7464) );
  CNR2X1 U8781 ( .A(n3848), .B(n6446), .Z(N833) );
  CEOX1 U8782 ( .A(N827), .B(mem_data1[809]), .Z(N7470) );
  CNR2X1 U8783 ( .A(n3848), .B(n6439), .Z(N827) );
  CEOX1 U8784 ( .A(N826), .B(mem_data1[808]), .Z(N7471) );
  CNR2X1 U8785 ( .A(n3841), .B(n6438), .Z(N826) );
  CEOX1 U8786 ( .A(N825), .B(mem_data1[807]), .Z(N7472) );
  CNR2X1 U8787 ( .A(n3840), .B(n6437), .Z(N825) );
  CEOX1 U8788 ( .A(N824), .B(mem_data1[806]), .Z(N7473) );
  CNR2X1 U8789 ( .A(n3839), .B(n6436), .Z(N824) );
  CEOX1 U8790 ( .A(N816), .B(mem_data1[798]), .Z(N7481) );
  CNR2X1 U8791 ( .A(n3835), .B(n6427), .Z(N816) );
  CEOX1 U8792 ( .A(N815), .B(mem_data1[797]), .Z(N7482) );
  CNR2X1 U8793 ( .A(n3834), .B(n6426), .Z(N815) );
  CEOX1 U8794 ( .A(N814), .B(mem_data1[796]), .Z(N7483) );
  CNR2X1 U8795 ( .A(n3853), .B(n6425), .Z(N814) );
  CEOX1 U8796 ( .A(N813), .B(mem_data1[795]), .Z(N7484) );
  CNR2X1 U8797 ( .A(n3852), .B(n6424), .Z(N813) );
  CEOX1 U8798 ( .A(N812), .B(mem_data1[794]), .Z(N7485) );
  CNR2X1 U8799 ( .A(n3851), .B(n6423), .Z(N812) );
  CEOX1 U8800 ( .A(N811), .B(mem_data1[793]), .Z(N7486) );
  CNR2X1 U8801 ( .A(n3850), .B(n6422), .Z(N811) );
  CEOX1 U8802 ( .A(N810), .B(mem_data1[792]), .Z(N7487) );
  CNR2X1 U8803 ( .A(n3849), .B(n6421), .Z(N810) );
  CEOX1 U8804 ( .A(N809), .B(mem_data1[791]), .Z(N7488) );
  CNR2X1 U8805 ( .A(n3848), .B(n6419), .Z(N809) );
  CEOX1 U8806 ( .A(N808), .B(mem_data1[790]), .Z(N7489) );
  CNR2X1 U8807 ( .A(n3847), .B(n6418), .Z(N808) );
  CEOX1 U8808 ( .A(N807), .B(mem_data1[789]), .Z(N7490) );
  CNR2X1 U8809 ( .A(n3846), .B(n6417), .Z(N807) );
  CEOX1 U8810 ( .A(N806), .B(mem_data1[788]), .Z(N7491) );
  CNR2X1 U8811 ( .A(n3845), .B(n6416), .Z(N806) );
  CEOX1 U8812 ( .A(N805), .B(mem_data1[787]), .Z(N7492) );
  CNR2X1 U8813 ( .A(n3844), .B(n6415), .Z(N805) );
  CEOX1 U8814 ( .A(N804), .B(mem_data1[786]), .Z(N7493) );
  CNR2X1 U8815 ( .A(n3836), .B(n6414), .Z(N804) );
  CEOX1 U8816 ( .A(N801), .B(mem_data1[783]), .Z(N7496) );
  CNR2X1 U8817 ( .A(n3834), .B(n6411), .Z(N801) );
  CEOX1 U8818 ( .A(N798), .B(mem_data1[780]), .Z(N7499) );
  CNR2X1 U8819 ( .A(n3842), .B(n6407), .Z(N798) );
  CEOX1 U8820 ( .A(N795), .B(mem_data1[777]), .Z(N7502) );
  CNR2X1 U8821 ( .A(n3838), .B(n6404), .Z(N795) );
  CEOX1 U8822 ( .A(N791), .B(mem_data1[773]), .Z(N7506) );
  CNR2X1 U8823 ( .A(n3834), .B(n6400), .Z(N791) );
  CEOX1 U8824 ( .A(N790), .B(mem_data1[772]), .Z(N7507) );
  CNR2X1 U8825 ( .A(n3846), .B(n6399), .Z(N790) );
  CEOX1 U8826 ( .A(N789), .B(mem_data1[771]), .Z(N7508) );
  CNR2X1 U8827 ( .A(n3853), .B(n6396), .Z(N789) );
  CEOX1 U8828 ( .A(N783), .B(mem_data1[765]), .Z(N7514) );
  CEOX1 U8829 ( .A(N782), .B(mem_data1[764]), .Z(N7515) );
  CEOX1 U8830 ( .A(N781), .B(mem_data1[763]), .Z(N7516) );
  CEOX1 U8831 ( .A(N780), .B(mem_data1[762]), .Z(N7517) );
  CEOX1 U8832 ( .A(N779), .B(mem_data1[761]), .Z(N7518) );
  CEOX1 U8833 ( .A(N778), .B(mem_data1[760]), .Z(N7519) );
  CEOX1 U8834 ( .A(N777), .B(mem_data1[759]), .Z(N7520) );
  CEOX1 U8835 ( .A(N776), .B(mem_data1[758]), .Z(N7521) );
  CEOX1 U8836 ( .A(N762), .B(mem_data1[744]), .Z(N7535) );
  CEOX1 U8837 ( .A(N758), .B(mem_data1[740]), .Z(N7539) );
  CEOX1 U8838 ( .A(N757), .B(mem_data1[739]), .Z(N7540) );
  CEOX1 U8839 ( .A(N756), .B(mem_data1[738]), .Z(N7541) );
  CEOX1 U8840 ( .A(N746), .B(mem_data1[728]), .Z(N7551) );
  CNR2X1 U8841 ( .A(n3832), .B(n6017), .Z(N746) );
  CEOX1 U8842 ( .A(N741), .B(mem_data1[723]), .Z(N7556) );
  CNR2X1 U8843 ( .A(n3825), .B(n6012), .Z(N741) );
  CEOX1 U8844 ( .A(N740), .B(mem_data1[722]), .Z(N7557) );
  CNR2X1 U8845 ( .A(n3826), .B(n6011), .Z(N740) );
  CEOX1 U8846 ( .A(N730), .B(mem_data1[712]), .Z(N7567) );
  CNR2X1 U8847 ( .A(n3823), .B(n6000), .Z(N730) );
  CEOX1 U8848 ( .A(N729), .B(mem_data1[711]), .Z(N7568) );
  CNR2X1 U8849 ( .A(n3819), .B(n5999), .Z(N729) );
  CEOX1 U8850 ( .A(N728), .B(mem_data1[710]), .Z(N7569) );
  CNR2X1 U8851 ( .A(n3820), .B(n5998), .Z(N728) );
  CEOX1 U8852 ( .A(N727), .B(mem_data1[709]), .Z(N7570) );
  CNR2X1 U8853 ( .A(n3815), .B(n5996), .Z(N727) );
  CEOX1 U8854 ( .A(N726), .B(mem_data1[708]), .Z(N7571) );
  CNR2X1 U8855 ( .A(n3816), .B(n5995), .Z(N726) );
  CEOX1 U8856 ( .A(N725), .B(mem_data1[707]), .Z(N7572) );
  CNR2X1 U8857 ( .A(n3817), .B(n5994), .Z(N725) );
  CEOX1 U8858 ( .A(N724), .B(mem_data1[706]), .Z(N7573) );
  CNR2X1 U8859 ( .A(n3832), .B(n5993), .Z(N724) );
  CEOX1 U8860 ( .A(N723), .B(mem_data1[705]), .Z(N7574) );
  CNR2X1 U8861 ( .A(n3833), .B(n5992), .Z(N723) );
  CEOX1 U8862 ( .A(N722), .B(mem_data1[704]), .Z(N7575) );
  CEOX1 U8863 ( .A(N721), .B(mem_data1[703]), .Z(N7576) );
  CNR2X1 U8864 ( .A(n3829), .B(n5990), .Z(N721) );
  CEOX1 U8865 ( .A(N720), .B(mem_data1[702]), .Z(N7577) );
  CNR2X1 U8866 ( .A(n3830), .B(n5989), .Z(N720) );
  CEOX1 U8867 ( .A(N719), .B(mem_data1[701]), .Z(N7578) );
  CNR2X1 U8868 ( .A(n3831), .B(n5988), .Z(N719) );
  CEOX1 U8869 ( .A(N718), .B(mem_data1[700]), .Z(N7579) );
  CNR2X1 U8870 ( .A(n3816), .B(n5987), .Z(N718) );
  CEOX1 U8871 ( .A(N717), .B(mem_data1[699]), .Z(N7580) );
  CNR2X1 U8872 ( .A(n3824), .B(n5984), .Z(N717) );
  CEOX1 U8873 ( .A(N716), .B(mem_data1[698]), .Z(N7581) );
  CNR2X1 U8874 ( .A(n3828), .B(n5983), .Z(N716) );
  CEOX1 U8875 ( .A(N715), .B(mem_data1[697]), .Z(N7582) );
  CNR2X1 U8876 ( .A(n3828), .B(n5982), .Z(N715) );
  CEOX1 U8877 ( .A(N714), .B(mem_data1[696]), .Z(N7583) );
  CNR2X1 U8878 ( .A(n3832), .B(n5981), .Z(N714) );
  CEOX1 U8879 ( .A(N713), .B(mem_data1[695]), .Z(N7584) );
  CNR2X1 U8880 ( .A(n3820), .B(n5980), .Z(N713) );
  CEOX1 U8881 ( .A(N712), .B(mem_data1[694]), .Z(N7585) );
  CNR2X1 U8882 ( .A(n3825), .B(n5979), .Z(N712) );
  CEOX1 U8883 ( .A(N711), .B(mem_data1[693]), .Z(N7586) );
  CNR2X1 U8884 ( .A(n3826), .B(n5978), .Z(N711) );
  CEOX1 U8885 ( .A(N710), .B(mem_data1[692]), .Z(N7587) );
  CNR2X1 U8886 ( .A(n3827), .B(n5977), .Z(N710) );
  CEOX1 U8887 ( .A(N706), .B(mem_data1[688]), .Z(N7591) );
  CNR2X1 U8888 ( .A(n3819), .B(n5972), .Z(N706) );
  CEOX1 U8889 ( .A(N705), .B(mem_data1[687]), .Z(N7592) );
  CNR2X1 U8890 ( .A(n3820), .B(n5971), .Z(N705) );
  CEOX1 U8891 ( .A(N704), .B(mem_data1[686]), .Z(N7593) );
  CNR2X1 U8892 ( .A(n3821), .B(n5970), .Z(N704) );
  CEOX1 U8893 ( .A(N698), .B(mem_data1[680]), .Z(N7599) );
  CNR2X1 U8894 ( .A(n3815), .B(n5964), .Z(N698) );
  CEOX1 U8895 ( .A(N693), .B(mem_data1[675]), .Z(N7604) );
  CNR2X1 U8896 ( .A(n3833), .B(n5958), .Z(N693) );
  CEOX1 U8897 ( .A(N692), .B(mem_data1[674]), .Z(N7605) );
  CNR2X1 U8898 ( .A(n3831), .B(n5957), .Z(N692) );
  CEOX1 U8899 ( .A(N688), .B(mem_data1[670]), .Z(N7609) );
  CNR2X1 U8900 ( .A(n3826), .B(n5953), .Z(N688) );
  CEOX1 U8901 ( .A(N685), .B(mem_data1[667]), .Z(N7612) );
  CNR2X1 U8902 ( .A(n3816), .B(n5949), .Z(N685) );
  CEOX1 U8903 ( .A(N678), .B(mem_data1[660]), .Z(N7619) );
  CNR2X1 U8904 ( .A(n3828), .B(n5942), .Z(N678) );
  CEOX1 U8905 ( .A(N677), .B(mem_data1[659]), .Z(N7620) );
  CNR2X1 U8906 ( .A(n3824), .B(n5940), .Z(N677) );
  CEOX1 U8907 ( .A(N676), .B(mem_data1[658]), .Z(N7621) );
  CNR2X1 U8908 ( .A(n3832), .B(n5939), .Z(N676) );
  CEOX1 U8909 ( .A(N666), .B(mem_data1[648]), .Z(N7631) );
  CNR2X1 U8910 ( .A(n3818), .B(n5928), .Z(N666) );
  CEOX1 U8911 ( .A(N665), .B(mem_data1[647]), .Z(N7632) );
  CNR2X1 U8912 ( .A(n3819), .B(n5927), .Z(N665) );
  CEOX1 U8913 ( .A(N664), .B(mem_data1[646]), .Z(N7633) );
  CNR2X1 U8914 ( .A(n3820), .B(n5926), .Z(N664) );
  CEOX1 U8915 ( .A(N660), .B(mem_data1[642]), .Z(N7637) );
  CNR2X1 U8916 ( .A(n3831), .B(n5922), .Z(N660) );
  CEOX1 U8917 ( .A(N659), .B(mem_data1[641]), .Z(N7638) );
  CNR2X1 U8918 ( .A(n3815), .B(n5921), .Z(N659) );
  CEOX1 U8919 ( .A(N658), .B(mem_data1[640]), .Z(N7639) );
  CEOX1 U8920 ( .A(N657), .B(mem_data1[639]), .Z(N7640) );
  CEOX1 U8921 ( .A(N656), .B(mem_data1[638]), .Z(N7641) );
  CEOX1 U8922 ( .A(N655), .B(mem_data1[637]), .Z(N7642) );
  CEOX1 U8923 ( .A(N654), .B(mem_data1[636]), .Z(N7643) );
  CEOX1 U8924 ( .A(N653), .B(mem_data1[635]), .Z(N7644) );
  CEOX1 U8925 ( .A(N652), .B(mem_data1[634]), .Z(N7645) );
  CEOX1 U8926 ( .A(N651), .B(mem_data1[633]), .Z(N7646) );
  CEOX1 U8927 ( .A(N650), .B(mem_data1[632]), .Z(N7647) );
  CEOX1 U8928 ( .A(N649), .B(mem_data1[631]), .Z(N7648) );
  CEOX1 U8929 ( .A(N648), .B(mem_data1[630]), .Z(N7649) );
  CEOX1 U8930 ( .A(N647), .B(mem_data1[629]), .Z(N7650) );
  CEOX1 U8931 ( .A(N646), .B(mem_data1[628]), .Z(N7651) );
  CEOX1 U8932 ( .A(N642), .B(mem_data1[624]), .Z(N7655) );
  CEOX1 U8933 ( .A(N641), .B(mem_data1[623]), .Z(N7656) );
  CEOX1 U8934 ( .A(N640), .B(mem_data1[622]), .Z(N7657) );
  CEOX1 U8935 ( .A(N634), .B(mem_data1[616]), .Z(N7663) );
  CEOX1 U8936 ( .A(N630), .B(mem_data1[612]), .Z(N7667) );
  CEOX1 U8937 ( .A(N629), .B(mem_data1[611]), .Z(N7668) );
  CEOX1 U8938 ( .A(N628), .B(mem_data1[610]), .Z(N7669) );
  CEOX1 U8939 ( .A(N618), .B(mem_data1[600]), .Z(N7679) );
  CNR2X1 U8940 ( .A(n3835), .B(n6017), .Z(N618) );
  CEOX1 U8941 ( .A(N613), .B(mem_data1[595]), .Z(N7684) );
  CNR2X1 U8942 ( .A(n3849), .B(n6012), .Z(N613) );
  CEOX1 U8943 ( .A(N612), .B(mem_data1[594]), .Z(N7685) );
  CNR2X1 U8944 ( .A(n3848), .B(n6011), .Z(N612) );
  CEOX1 U8945 ( .A(N602), .B(mem_data1[584]), .Z(N7695) );
  CNR2X1 U8946 ( .A(n3845), .B(n6000), .Z(N602) );
  CEOX1 U8947 ( .A(N601), .B(mem_data1[583]), .Z(N7696) );
  CNR2X1 U8948 ( .A(n3847), .B(n5999), .Z(N601) );
  CEOX1 U8949 ( .A(N600), .B(mem_data1[582]), .Z(N7697) );
  CNR2X1 U8950 ( .A(n3841), .B(n5998), .Z(N600) );
  CEOX1 U8951 ( .A(N599), .B(mem_data1[581]), .Z(N7698) );
  CNR2X1 U8952 ( .A(n3840), .B(n5996), .Z(N599) );
  CEOX1 U8953 ( .A(N598), .B(mem_data1[580]), .Z(N7699) );
  CNR2X1 U8954 ( .A(n3839), .B(n5995), .Z(N598) );
  CEOX1 U8955 ( .A(N597), .B(mem_data1[579]), .Z(N7700) );
  CNR2X1 U8956 ( .A(n3837), .B(n5994), .Z(N597) );
  CEOX1 U8957 ( .A(N596), .B(mem_data1[578]), .Z(N7701) );
  CNR2X1 U8958 ( .A(n3836), .B(n5993), .Z(N596) );
  CEOX1 U8959 ( .A(N592), .B(mem_data1[574]), .Z(N7705) );
  CNR2X1 U8960 ( .A(n3852), .B(n5989), .Z(N592) );
  CEOX1 U8961 ( .A(N591), .B(mem_data1[573]), .Z(N7706) );
  CNR2X1 U8962 ( .A(n3843), .B(n5988), .Z(N591) );
  CEOX1 U8963 ( .A(N590), .B(mem_data1[572]), .Z(N7707) );
  CNR2X1 U8964 ( .A(n3851), .B(n5987), .Z(N590) );
  CEOX1 U8965 ( .A(N589), .B(mem_data1[571]), .Z(N7708) );
  CNR2X1 U8966 ( .A(n3850), .B(n5984), .Z(N589) );
  CEOX1 U8967 ( .A(N588), .B(mem_data1[570]), .Z(N7709) );
  CNR2X1 U8968 ( .A(n3849), .B(n5983), .Z(N588) );
  CEOX1 U8969 ( .A(N587), .B(mem_data1[569]), .Z(N7710) );
  CNR2X1 U8970 ( .A(n3844), .B(n5982), .Z(N587) );
  CEOX1 U8971 ( .A(N586), .B(mem_data1[568]), .Z(N7711) );
  CNR2X1 U8972 ( .A(n3846), .B(n5981), .Z(N586) );
  CEOX1 U8973 ( .A(N585), .B(mem_data1[567]), .Z(N7712) );
  CNR2X1 U8974 ( .A(n3843), .B(n5980), .Z(N585) );
  CEOX1 U8975 ( .A(N584), .B(mem_data1[566]), .Z(N7713) );
  CNR2X1 U8976 ( .A(n3842), .B(n5979), .Z(N584) );
  CEOX1 U8977 ( .A(N583), .B(mem_data1[565]), .Z(N7714) );
  CNR2X1 U8978 ( .A(n3846), .B(n5978), .Z(N583) );
  CEOX1 U8979 ( .A(N582), .B(mem_data1[564]), .Z(N7715) );
  CNR2X1 U8980 ( .A(n3847), .B(n5977), .Z(N582) );
  CEOX1 U8981 ( .A(N578), .B(mem_data1[560]), .Z(N7719) );
  CNR2X1 U8982 ( .A(n3843), .B(n5972), .Z(N578) );
  CEOX1 U8983 ( .A(N577), .B(mem_data1[559]), .Z(N7720) );
  CNR2X1 U8984 ( .A(n3841), .B(n5971), .Z(N577) );
  CEOX1 U8985 ( .A(N576), .B(mem_data1[558]), .Z(N7721) );
  CNR2X1 U8986 ( .A(n3840), .B(n5970), .Z(N576) );
  CEOX1 U8987 ( .A(N570), .B(mem_data1[552]), .Z(N7727) );
  CNR2X1 U8988 ( .A(n3835), .B(n5964), .Z(N570) );
  CEOX1 U8989 ( .A(N566), .B(mem_data1[548]), .Z(N7731) );
  CNR2X1 U8990 ( .A(n3839), .B(n5959), .Z(N566) );
  CEOX1 U8991 ( .A(N565), .B(mem_data1[547]), .Z(N7732) );
  CNR2X1 U8992 ( .A(n3845), .B(n5958), .Z(N565) );
  CEOX1 U8993 ( .A(N564), .B(mem_data1[546]), .Z(N7733) );
  CNR2X1 U8994 ( .A(n3853), .B(n5957), .Z(N564) );
  CEOX1 U8995 ( .A(N560), .B(mem_data1[542]), .Z(N7737) );
  CNR2X1 U8996 ( .A(n3849), .B(n5953), .Z(N560) );
  CEOX1 U8997 ( .A(N557), .B(mem_data1[539]), .Z(N7740) );
  CNR2X1 U8998 ( .A(n3845), .B(n5949), .Z(N557) );
  CEOX1 U8999 ( .A(N550), .B(mem_data1[532]), .Z(N7747) );
  CNR2X1 U9000 ( .A(n3838), .B(n5942), .Z(N550) );
  CEOX1 U9001 ( .A(N549), .B(mem_data1[531]), .Z(N7748) );
  CNR2X1 U9002 ( .A(n3844), .B(n5940), .Z(N549) );
  CEOX1 U9003 ( .A(N548), .B(mem_data1[530]), .Z(N7749) );
  CNR2X1 U9004 ( .A(n3837), .B(n5939), .Z(N548) );
  CEOX1 U9005 ( .A(N538), .B(mem_data1[520]), .Z(N7759) );
  CNR2X1 U9006 ( .A(n3851), .B(n5928), .Z(N538) );
  CEOX1 U9007 ( .A(N537), .B(mem_data1[519]), .Z(N7760) );
  CNR2X1 U9008 ( .A(n3840), .B(n5927), .Z(N537) );
  CEOX1 U9009 ( .A(N536), .B(mem_data1[518]), .Z(N7761) );
  CNR2X1 U9010 ( .A(n3849), .B(n5926), .Z(N536) );
  CEOX1 U9011 ( .A(N532), .B(mem_data1[514]), .Z(N7765) );
  CNR2X1 U9012 ( .A(n3835), .B(n5922), .Z(N532) );
  CEOX1 U9013 ( .A(N528), .B(mem_data1[510]), .Z(N7769) );
  CEOX1 U9014 ( .A(N527), .B(mem_data1[509]), .Z(N7770) );
  CEOX1 U9015 ( .A(N526), .B(mem_data1[508]), .Z(N7771) );
  CEOX1 U9016 ( .A(N525), .B(mem_data1[507]), .Z(N7772) );
  CEOX1 U9017 ( .A(N524), .B(mem_data1[506]), .Z(N7773) );
  CEOX1 U9018 ( .A(N519), .B(mem_data1[501]), .Z(N7778) );
  CEOX1 U9019 ( .A(N493), .B(mem_data1[475]), .Z(N7804) );
  CNR2X1 U9020 ( .A(n3833), .B(n5457), .Z(N493) );
  CEOX1 U9021 ( .A(N492), .B(mem_data1[474]), .Z(N7805) );
  CNR2X1 U9022 ( .A(n3828), .B(n5456), .Z(N492) );
  CEOX1 U9023 ( .A(N491), .B(mem_data1[473]), .Z(N7806) );
  CNR2X1 U9024 ( .A(n3829), .B(n5455), .Z(N491) );
  CEOX1 U9025 ( .A(N490), .B(mem_data1[472]), .Z(N7807) );
  CNR2X1 U9026 ( .A(n3830), .B(n5454), .Z(N490) );
  CEOX1 U9027 ( .A(N489), .B(mem_data1[471]), .Z(N7808) );
  CNR2X1 U9028 ( .A(n3825), .B(n5453), .Z(N489) );
  CEOX1 U9029 ( .A(N488), .B(mem_data1[470]), .Z(N7809) );
  CNR2X1 U9030 ( .A(n3826), .B(n5452), .Z(N488) );
  CEOX1 U9031 ( .A(N487), .B(mem_data1[469]), .Z(N7810) );
  CNR2X1 U9032 ( .A(n3827), .B(n5450), .Z(N487) );
  CEOX1 U9033 ( .A(N486), .B(mem_data1[468]), .Z(N7811) );
  CNR2X1 U9034 ( .A(n3822), .B(n5449), .Z(N486) );
  CEOX1 U9035 ( .A(N485), .B(mem_data1[467]), .Z(N7812) );
  CNR2IX1 U9036 ( .B(n3841), .A(n5448), .Z(N485) );
  CEOX1 U9037 ( .A(N479), .B(mem_data1[461]), .Z(N7818) );
  CNR2X1 U9038 ( .A(n3817), .B(n5442), .Z(N479) );
  CEOX1 U9039 ( .A(N478), .B(mem_data1[460]), .Z(N7819) );
  CNR2X1 U9040 ( .A(n3816), .B(n5441), .Z(N478) );
  CEOX1 U9041 ( .A(N477), .B(mem_data1[459]), .Z(N7820) );
  CNR2IX1 U9042 ( .B(n3847), .A(n5439), .Z(N477) );
  CEOX1 U9043 ( .A(N476), .B(mem_data1[458]), .Z(N7821) );
  CNR2X1 U9044 ( .A(n3833), .B(n5438), .Z(N476) );
  CEOX1 U9045 ( .A(N475), .B(mem_data1[457]), .Z(N7822) );
  CNR2X1 U9046 ( .A(n3828), .B(n5437), .Z(N475) );
  CEOX1 U9047 ( .A(N469), .B(mem_data1[451]), .Z(N7828) );
  CNR2X1 U9048 ( .A(n3828), .B(n5431), .Z(N469) );
  CEOX1 U9049 ( .A(N468), .B(mem_data1[450]), .Z(N7829) );
  CNR2X1 U9050 ( .A(n3823), .B(n5430), .Z(N468) );
  CEOX1 U9051 ( .A(N467), .B(mem_data1[449]), .Z(N7830) );
  CNR2X1 U9052 ( .A(n3824), .B(n5428), .Z(N467) );
  CEOX1 U9053 ( .A(N429), .B(mem_data1[411]), .Z(N7868) );
  CNR2X1 U9054 ( .A(n3815), .B(n5387), .Z(N429) );
  CEOX1 U9055 ( .A(N428), .B(mem_data1[410]), .Z(N7869) );
  CNR2X1 U9056 ( .A(n3819), .B(n5386), .Z(N428) );
  CEOX1 U9057 ( .A(N427), .B(mem_data1[409]), .Z(N7870) );
  CNR2X1 U9058 ( .A(n3832), .B(n5384), .Z(N427) );
  CEOX1 U9059 ( .A(N426), .B(mem_data1[408]), .Z(N7871) );
  CNR2X1 U9060 ( .A(n3833), .B(n5383), .Z(N426) );
  CEOX1 U9061 ( .A(N425), .B(mem_data1[407]), .Z(N7872) );
  CNR2X1 U9062 ( .A(n3814), .B(n5382), .Z(N425) );
  CEOX1 U9063 ( .A(N424), .B(mem_data1[406]), .Z(N7873) );
  CNR2X1 U9064 ( .A(n3829), .B(n5381), .Z(N424) );
  CEOX1 U9065 ( .A(N423), .B(mem_data1[405]), .Z(N7874) );
  CNR2X1 U9066 ( .A(n3830), .B(n5380), .Z(N423) );
  CEOX1 U9067 ( .A(N415), .B(mem_data1[397]), .Z(N7882) );
  CNR2X1 U9068 ( .A(n3816), .B(n5370), .Z(N415) );
  CEOX1 U9069 ( .A(N411), .B(mem_data1[393]), .Z(N7886) );
  CNR2X1 U9070 ( .A(n3824), .B(n5366), .Z(N411) );
  CEOX1 U9071 ( .A(N407), .B(mem_data1[389]), .Z(N7890) );
  CNR2IX1 U9072 ( .B(n3842), .A(n5361), .Z(N407) );
  CEOX1 U9073 ( .A(N406), .B(mem_data1[388]), .Z(N7891) );
  CNR2X1 U9074 ( .A(n3819), .B(n5360), .Z(N406) );
  CEOX1 U9075 ( .A(N405), .B(mem_data1[387]), .Z(N7892) );
  CNR2X1 U9076 ( .A(n3830), .B(n5359), .Z(N405) );
  CEOX1 U9077 ( .A(N404), .B(mem_data1[386]), .Z(N7893) );
  CNR2X1 U9078 ( .A(n3820), .B(n5358), .Z(N404) );
  CEOX1 U9079 ( .A(N403), .B(mem_data1[385]), .Z(N7894) );
  CNR2X1 U9080 ( .A(n3821), .B(n5357), .Z(N403) );
  CEOX1 U9081 ( .A(N364), .B(mem_data1[346]), .Z(N7933) );
  CNR2X1 U9082 ( .A(n3850), .B(n5456), .Z(N364) );
  CEOX1 U9083 ( .A(N363), .B(mem_data1[345]), .Z(N7934) );
  CNR2X1 U9084 ( .A(n3849), .B(n5455), .Z(N363) );
  CEOX1 U9085 ( .A(N362), .B(mem_data1[344]), .Z(N7935) );
  CNR2X1 U9086 ( .A(n3848), .B(n5454), .Z(N362) );
  CEOX1 U9087 ( .A(N361), .B(mem_data1[343]), .Z(N7936) );
  CNR2X1 U9088 ( .A(n3847), .B(n5453), .Z(N361) );
  CEOX1 U9089 ( .A(N360), .B(mem_data1[342]), .Z(N7937) );
  CNR2X1 U9090 ( .A(n3846), .B(n5452), .Z(N360) );
  CEOX1 U9091 ( .A(N359), .B(mem_data1[341]), .Z(N7938) );
  CNR2X1 U9092 ( .A(n3845), .B(n5450), .Z(N359) );
  CEOX1 U9093 ( .A(mem_data1[337]), .B(N355), .Z(N7942) );
  CNR2IX1 U9094 ( .B(n3815), .A(n5446), .Z(N355) );
  CEOX1 U9095 ( .A(N351), .B(mem_data1[333]), .Z(N7946) );
  CNR2X1 U9096 ( .A(n3849), .B(n5442), .Z(N351) );
  CEOX1 U9097 ( .A(N347), .B(mem_data1[329]), .Z(N7950) );
  CNR2X1 U9098 ( .A(n3837), .B(n5437), .Z(N347) );
  CEOX1 U9099 ( .A(N341), .B(mem_data1[323]), .Z(N7956) );
  CNR2X1 U9100 ( .A(n3851), .B(n5431), .Z(N341) );
  CEOX1 U9101 ( .A(N340), .B(mem_data1[322]), .Z(N7957) );
  CNR2X1 U9102 ( .A(n3850), .B(n5430), .Z(N340) );
  CEOX1 U9103 ( .A(N339), .B(mem_data1[321]), .Z(N7958) );
  CNR2X1 U9104 ( .A(n3849), .B(n5428), .Z(N339) );
  CEOX1 U9105 ( .A(N301), .B(mem_data1[283]), .Z(N7996) );
  CNR2X1 U9106 ( .A(n3835), .B(n5387), .Z(N301) );
  CEOX1 U9107 ( .A(N300), .B(mem_data1[282]), .Z(N7997) );
  CNR2X1 U9108 ( .A(n3839), .B(n5386), .Z(N300) );
  CEOX1 U9109 ( .A(N299), .B(mem_data1[281]), .Z(N7998) );
  CNR2X1 U9110 ( .A(n3838), .B(n5384), .Z(N299) );
  CEOX1 U9111 ( .A(N298), .B(mem_data1[280]), .Z(N7999) );
  CNR2X1 U9112 ( .A(n3837), .B(n5383), .Z(N298) );
  CEOX1 U9113 ( .A(N297), .B(mem_data1[279]), .Z(N8000) );
  CNR2X1 U9114 ( .A(n3840), .B(n5382), .Z(N297) );
  CEOX1 U9115 ( .A(N296), .B(mem_data1[278]), .Z(N8001) );
  CNR2X1 U9116 ( .A(n3838), .B(n5381), .Z(N296) );
  CEOX1 U9117 ( .A(N295), .B(mem_data1[277]), .Z(N8002) );
  CNR2X1 U9118 ( .A(n3839), .B(n5380), .Z(N295) );
  CEOX1 U9119 ( .A(N291), .B(mem_data1[273]), .Z(N8006) );
  CNR2IX1 U9120 ( .B(n3816), .A(n5376), .Z(N291) );
  CEOX1 U9121 ( .A(N288), .B(mem_data1[270]), .Z(N8009) );
  CNR2X1 U9122 ( .A(n3851), .B(n5371), .Z(N288) );
  CEOX1 U9123 ( .A(N287), .B(mem_data1[269]), .Z(N8010) );
  CNR2X1 U9124 ( .A(n3849), .B(n5370), .Z(N287) );
  CEOX1 U9125 ( .A(N283), .B(mem_data1[265]), .Z(N8014) );
  CNR2X1 U9126 ( .A(n3834), .B(n5366), .Z(N283) );
  CEOX1 U9127 ( .A(N277), .B(mem_data1[259]), .Z(N8020) );
  CNR2X1 U9128 ( .A(n3836), .B(n5359), .Z(N277) );
  CEOX1 U9129 ( .A(N276), .B(mem_data1[258]), .Z(N8021) );
  CNR2X1 U9130 ( .A(n3835), .B(n5358), .Z(N276) );
  CEOX1 U9131 ( .A(N275), .B(mem_data1[257]), .Z(N8022) );
  CNR2X1 U9132 ( .A(n3837), .B(n5357), .Z(N275) );
  CEOX1 U9133 ( .A(N254), .B(mem_data1[236]), .Z(N8043) );
  CEOX1 U9134 ( .A(N253), .B(mem_data1[235]), .Z(N8044) );
  CEOX1 U9135 ( .A(N252), .B(mem_data1[234]), .Z(N8045) );
  CEOX1 U9136 ( .A(N243), .B(mem_data1[225]), .Z(N8054) );
  CEOX1 U9137 ( .A(N242), .B(mem_data1[224]), .Z(N8055) );
  CNR2X1 U9138 ( .A(n3818), .B(n6475), .Z(N242) );
  CEOX1 U9139 ( .A(N241), .B(mem_data1[223]), .Z(N8056) );
  CNR2X1 U9140 ( .A(n3822), .B(n6464), .Z(N241) );
  CEOX1 U9141 ( .A(N238), .B(mem_data1[220]), .Z(N8059) );
  CNR2X1 U9142 ( .A(n3823), .B(n6431), .Z(N238) );
  CEOX1 U9143 ( .A(N237), .B(mem_data1[219]), .Z(N8060) );
  CNR2X1 U9144 ( .A(n3815), .B(n6420), .Z(N237) );
  CEOX1 U9145 ( .A(N236), .B(mem_data1[218]), .Z(N8061) );
  CNR2X1 U9146 ( .A(n3816), .B(n6409), .Z(N236) );
  CEOX1 U9147 ( .A(N235), .B(mem_data1[217]), .Z(N8062) );
  CNR2X1 U9148 ( .A(n3817), .B(n6397), .Z(N235) );
  CEOX1 U9149 ( .A(N234), .B(mem_data1[216]), .Z(N8063) );
  CNR2X1 U9150 ( .A(n3832), .B(n6380), .Z(N234) );
  CEOX1 U9151 ( .A(N233), .B(mem_data1[215]), .Z(N8064) );
  CNR2X1 U9152 ( .A(n3833), .B(n6359), .Z(N233) );
  CEOX1 U9153 ( .A(N232), .B(mem_data1[214]), .Z(N8065) );
  CNR2X1 U9154 ( .A(n3822), .B(n6338), .Z(N232) );
  CEOX1 U9155 ( .A(N231), .B(mem_data1[213]), .Z(N8066) );
  CNR2X1 U9156 ( .A(n3829), .B(n6322), .Z(N231) );
  CEOX1 U9157 ( .A(N230), .B(mem_data1[212]), .Z(N8067) );
  CNR2X1 U9158 ( .A(n3830), .B(n6311), .Z(N230) );
  CEOX1 U9159 ( .A(N229), .B(mem_data1[211]), .Z(N8068) );
  CNR2X1 U9160 ( .A(n3831), .B(n6300), .Z(N229) );
  CEOX1 U9161 ( .A(N228), .B(mem_data1[210]), .Z(N8069) );
  CNR2X1 U9162 ( .A(n3826), .B(n6287), .Z(N228) );
  CEOX1 U9163 ( .A(N227), .B(mem_data1[209]), .Z(N8070) );
  CNR2X1 U9164 ( .A(n3827), .B(n6266), .Z(N227) );
  CEOX1 U9165 ( .A(N226), .B(mem_data1[208]), .Z(N8071) );
  CNR2X1 U9166 ( .A(n3828), .B(n6245), .Z(N226) );
  CEOX1 U9167 ( .A(N225), .B(mem_data1[207]), .Z(N8072) );
  CNR2X1 U9168 ( .A(n3821), .B(n6224), .Z(N225) );
  CEOX1 U9169 ( .A(N224), .B(mem_data1[206]), .Z(N8073) );
  CNR2X1 U9170 ( .A(n3824), .B(n6203), .Z(N224) );
  CEOX1 U9171 ( .A(N223), .B(mem_data1[205]), .Z(N8074) );
  CNR2X1 U9172 ( .A(n3825), .B(n6182), .Z(N223) );
  CEOX1 U9173 ( .A(N222), .B(mem_data1[204]), .Z(N8075) );
  CNR2X1 U9174 ( .A(n3833), .B(n6155), .Z(N222) );
  CEOX1 U9175 ( .A(N221), .B(mem_data1[203]), .Z(N8076) );
  CNR2X1 U9176 ( .A(n3829), .B(n6125), .Z(N221) );
  CEOX1 U9177 ( .A(N220), .B(mem_data1[202]), .Z(N8077) );
  CNR2X1 U9178 ( .A(n3817), .B(n6085), .Z(N220) );
  CEOX1 U9179 ( .A(N219), .B(mem_data1[201]), .Z(N8078) );
  CNR2X1 U9180 ( .A(n3822), .B(n6036), .Z(N219) );
  CEOX1 U9181 ( .A(N218), .B(mem_data1[200]), .Z(N8079) );
  CNR2X1 U9182 ( .A(n3823), .B(n6019), .Z(N218) );
  CEOX1 U9183 ( .A(N217), .B(mem_data1[199]), .Z(N8080) );
  CNR2X1 U9184 ( .A(n3825), .B(n6008), .Z(N217) );
  CEOX1 U9185 ( .A(N216), .B(mem_data1[198]), .Z(N8081) );
  CNR2X1 U9186 ( .A(n3819), .B(n5997), .Z(N216) );
  CEOX1 U9187 ( .A(N215), .B(mem_data1[197]), .Z(N8082) );
  CNR2X1 U9188 ( .A(n3820), .B(n5985), .Z(N215) );
  CEOX1 U9189 ( .A(N214), .B(mem_data1[196]), .Z(N8083) );
  CNR2X1 U9190 ( .A(n3821), .B(n5974), .Z(N214) );
  CEOX1 U9191 ( .A(N213), .B(mem_data1[195]), .Z(N8084) );
  CNR2X1 U9192 ( .A(n3816), .B(n5963), .Z(N213) );
  CEOX1 U9193 ( .A(N212), .B(mem_data1[194]), .Z(N8085) );
  CNR2X1 U9194 ( .A(n3817), .B(n5952), .Z(N212) );
  CEOX1 U9195 ( .A(N211), .B(mem_data1[193]), .Z(N8086) );
  CNR2X1 U9196 ( .A(n3818), .B(n5941), .Z(N211) );
  CEOX1 U9197 ( .A(N210), .B(mem_data1[192]), .Z(N8087) );
  CNR2X1 U9198 ( .A(n3833), .B(n5930), .Z(N210) );
  CEOX1 U9199 ( .A(N209), .B(mem_data1[191]), .Z(N8088) );
  CNR2X1 U9200 ( .A(n3829), .B(n5919), .Z(N209) );
  CEOX1 U9201 ( .A(N205), .B(mem_data1[187]), .Z(N8092) );
  CNR2X1 U9202 ( .A(n3832), .B(n5843), .Z(N205) );
  CEOX1 U9203 ( .A(N204), .B(mem_data1[186]), .Z(N8093) );
  CNR2X1 U9204 ( .A(n3816), .B(n5832), .Z(N204) );
  CEOX1 U9205 ( .A(N203), .B(mem_data1[185]), .Z(N8094) );
  CNR2X1 U9206 ( .A(n3820), .B(n5821), .Z(N203) );
  CEOX1 U9207 ( .A(N202), .B(mem_data1[184]), .Z(N8095) );
  CNR2X1 U9208 ( .A(n3829), .B(n5804), .Z(N202) );
  CEOX1 U9209 ( .A(N201), .B(mem_data1[183]), .Z(N8096) );
  CNR2X1 U9210 ( .A(n3824), .B(n5783), .Z(N201) );
  CEOX1 U9211 ( .A(N200), .B(mem_data1[182]), .Z(N8097) );
  CNR2X1 U9212 ( .A(n3832), .B(n5762), .Z(N200) );
  CEOX1 U9213 ( .A(N199), .B(mem_data1[181]), .Z(N8098) );
  CNR2X1 U9214 ( .A(n3828), .B(n5742), .Z(N199) );
  CEOX1 U9215 ( .A(N198), .B(mem_data1[180]), .Z(N8099) );
  CNR2X1 U9216 ( .A(n3826), .B(n5721), .Z(N198) );
  CEOX1 U9217 ( .A(N197), .B(mem_data1[179]), .Z(N8100) );
  CNR2X1 U9218 ( .A(n3827), .B(n5692), .Z(N197) );
  CEOX1 U9219 ( .A(N196), .B(mem_data1[178]), .Z(N8101) );
  CNR2X1 U9220 ( .A(n3828), .B(n5639), .Z(N196) );
  CEOX1 U9221 ( .A(N195), .B(mem_data1[177]), .Z(N8102) );
  CNR2X1 U9222 ( .A(n3823), .B(n5567), .Z(N195) );
  CEOX1 U9223 ( .A(N194), .B(mem_data1[176]), .Z(N8103) );
  CEOX1 U9224 ( .A(N193), .B(mem_data1[175]), .Z(N8104) );
  CNR2X1 U9225 ( .A(n3825), .B(n5462), .Z(N193) );
  CEOX1 U9226 ( .A(N191), .B(mem_data1[173]), .Z(N8106) );
  CNR2X1 U9227 ( .A(n3821), .B(n5440), .Z(N191) );
  CEOX1 U9228 ( .A(N190), .B(mem_data1[172]), .Z(N8107) );
  CNR2X1 U9229 ( .A(n3822), .B(n5429), .Z(N190) );
  CEOX1 U9230 ( .A(N189), .B(mem_data1[171]), .Z(N8108) );
  CNR2X1 U9231 ( .A(n3817), .B(n5418), .Z(N189) );
  CEOX1 U9232 ( .A(N188), .B(mem_data1[170]), .Z(N8109) );
  CNR2X1 U9233 ( .A(n3818), .B(n5407), .Z(N188) );
  CEOX1 U9234 ( .A(N187), .B(mem_data1[169]), .Z(N8110) );
  CNR2X1 U9235 ( .A(n3819), .B(n5396), .Z(N187) );
  CEOX1 U9236 ( .A(N186), .B(mem_data1[168]), .Z(N8111) );
  CNR2X1 U9237 ( .A(n3832), .B(n5385), .Z(N186) );
  CEOX1 U9238 ( .A(N185), .B(mem_data1[167]), .Z(N8112) );
  CNR2X1 U9239 ( .A(n3815), .B(n5373), .Z(N185) );
  CEOX1 U9240 ( .A(N184), .B(mem_data1[166]), .Z(N8113) );
  CNR2X1 U9241 ( .A(n3827), .B(n5362), .Z(N184) );
  CEOX1 U9242 ( .A(N183), .B(mem_data1[165]), .Z(N8114) );
  CNR2X1 U9243 ( .A(n3815), .B(n5347), .Z(N183) );
  CEOX1 U9244 ( .A(N179), .B(mem_data1[161]), .Z(N8118) );
  CNR2X1 U9245 ( .A(n3831), .B(n5276), .Z(N179) );
  CEOX1 U9246 ( .A(N178), .B(mem_data1[160]), .Z(N8119) );
  CNR2X1 U9247 ( .A(n3830), .B(n5265), .Z(N178) );
  CEOX1 U9248 ( .A(N177), .B(mem_data1[159]), .Z(N8120) );
  CNR2X1 U9249 ( .A(n3831), .B(n5254), .Z(N177) );
  CEOX1 U9250 ( .A(N175), .B(mem_data1[157]), .Z(N8122) );
  CNR2X1 U9251 ( .A(n3827), .B(n5211), .Z(N175) );
  CEOX1 U9252 ( .A(N174), .B(mem_data1[156]), .Z(N8123) );
  CNR2X1 U9253 ( .A(n3828), .B(n5190), .Z(N174) );
  CEOX1 U9254 ( .A(N172), .B(mem_data1[154]), .Z(N8125) );
  CNR2X1 U9255 ( .A(n3824), .B(n5147), .Z(N172) );
  CEOX1 U9256 ( .A(N171), .B(mem_data1[153]), .Z(N8126) );
  CNR2X1 U9257 ( .A(n3825), .B(n5112), .Z(N171) );
  CEOX1 U9258 ( .A(N170), .B(mem_data1[152]), .Z(N8127) );
  CNR2X1 U9259 ( .A(n3826), .B(n5047), .Z(N170) );
  CEOX1 U9260 ( .A(N169), .B(mem_data1[151]), .Z(N8128) );
  CNR2X1 U9261 ( .A(n3821), .B(n4977), .Z(N169) );
  CEOX1 U9262 ( .A(N168), .B(mem_data1[150]), .Z(N8129) );
  CNR2X1 U9263 ( .A(n3822), .B(n4922), .Z(N168) );
  CEOX1 U9264 ( .A(N167), .B(mem_data1[149]), .Z(N8130) );
  CNR2X1 U9265 ( .A(n3823), .B(n4903), .Z(N167) );
  CEOX1 U9266 ( .A(N166), .B(mem_data1[148]), .Z(N8131) );
  CNR2X1 U9267 ( .A(n3818), .B(n4892), .Z(N166) );
  CEOX1 U9268 ( .A(N165), .B(mem_data1[147]), .Z(N8132) );
  CNR2X1 U9269 ( .A(n3819), .B(n4880), .Z(N165) );
  CEOX1 U9270 ( .A(N164), .B(mem_data1[146]), .Z(N8133) );
  CNR2X1 U9271 ( .A(n3820), .B(n4867), .Z(N164) );
  CEOX1 U9272 ( .A(N163), .B(mem_data1[145]), .Z(N8134) );
  CNR2X1 U9273 ( .A(n3830), .B(n4846), .Z(N163) );
  CEOX1 U9274 ( .A(N162), .B(mem_data1[144]), .Z(N8135) );
  CNR2X1 U9275 ( .A(n3826), .B(n4825), .Z(N162) );
  CEOX1 U9276 ( .A(N161), .B(mem_data1[143]), .Z(N8136) );
  CNR2X1 U9277 ( .A(n3833), .B(n4805), .Z(N161) );
  CEOX1 U9278 ( .A(N160), .B(mem_data1[142]), .Z(N8137) );
  CEOX1 U9279 ( .A(N159), .B(mem_data1[141]), .Z(N8138) );
  CEOX1 U9280 ( .A(N158), .B(mem_data1[140]), .Z(N8139) );
  CEOX1 U9281 ( .A(N157), .B(mem_data1[139]), .Z(N8140) );
  CEOX1 U9282 ( .A(N156), .B(mem_data1[138]), .Z(N8141) );
  CEOX1 U9283 ( .A(N155), .B(mem_data1[137]), .Z(N8142) );
  CEOX1 U9284 ( .A(N154), .B(mem_data1[136]), .Z(N8143) );
  CNR2X1 U9285 ( .A(n3831), .B(n6398), .Z(N154) );
  CEOX1 U9286 ( .A(N153), .B(mem_data1[135]), .Z(N8144) );
  CNR2X1 U9287 ( .A(n3832), .B(n6225), .Z(N153) );
  CEOX1 U9288 ( .A(N152), .B(mem_data1[134]), .Z(N8145) );
  CNR2X1 U9289 ( .A(n3833), .B(n5986), .Z(N152) );
  CEOX1 U9290 ( .A(N151), .B(mem_data1[133]), .Z(N8146) );
  CNR2X1 U9291 ( .A(n3828), .B(n5844), .Z(N151) );
  CEOX1 U9292 ( .A(N149), .B(mem_data1[131]), .Z(N8148) );
  CNR2X1 U9293 ( .A(n3830), .B(n5374), .Z(N149) );
  CEOX1 U9294 ( .A(N148), .B(mem_data1[130]), .Z(N8149) );
  CNR2X1 U9295 ( .A(n3825), .B(n5212), .Z(N148) );
  CEOX1 U9296 ( .A(N147), .B(mem_data1[129]), .Z(N8150) );
  CNR2X1 U9297 ( .A(n3826), .B(n4881), .Z(N147) );
  CEOX1 U9298 ( .A(N131), .B(mem_data1[113]), .Z(N8166) );
  CEOX1 U9299 ( .A(N130), .B(mem_data1[112]), .Z(N8167) );
  CEOX1 U9300 ( .A(N125), .B(mem_data1[107]), .Z(N8172) );
  CEOX1 U9301 ( .A(N124), .B(mem_data1[106]), .Z(N8173) );
  CND2X1 U9302 ( .A(n4827), .B(n3729), .Z(n4631) );
  CEOX1 U9303 ( .A(N110), .B(mem_data1[92]), .Z(N8187) );
  CNR2X1 U9304 ( .A(n3836), .B(n6431), .Z(N110) );
  CEOX1 U9305 ( .A(N109), .B(mem_data1[91]), .Z(N8188) );
  CNR2X1 U9306 ( .A(n3836), .B(n6420), .Z(N109) );
  CEOX1 U9307 ( .A(N108), .B(mem_data1[90]), .Z(N8189) );
  CNR2X1 U9308 ( .A(n3835), .B(n6409), .Z(N108) );
  CEOX1 U9309 ( .A(N107), .B(mem_data1[89]), .Z(N8190) );
  CNR2X1 U9310 ( .A(n3848), .B(n6397), .Z(N107) );
  CEOX1 U9311 ( .A(N106), .B(mem_data1[88]), .Z(N8191) );
  CNR2X1 U9312 ( .A(n3847), .B(n6380), .Z(N106) );
  CEOX1 U9313 ( .A(N105), .B(mem_data1[87]), .Z(N8192) );
  CNR2X1 U9314 ( .A(n3846), .B(n6359), .Z(N105) );
  CEOX1 U9315 ( .A(N104), .B(mem_data1[86]), .Z(N8193) );
  CNR2X1 U9316 ( .A(n3845), .B(n6338), .Z(N104) );
  CEOX1 U9317 ( .A(N103), .B(mem_data1[85]), .Z(N8194) );
  CNR2X1 U9318 ( .A(n3840), .B(n6322), .Z(N103) );
  CEOX1 U9319 ( .A(N102), .B(mem_data1[84]), .Z(N8195) );
  CNR2X1 U9320 ( .A(n3834), .B(n6311), .Z(N102) );
  CEOX1 U9321 ( .A(N101), .B(mem_data1[83]), .Z(N8196) );
  CNR2X1 U9322 ( .A(n3853), .B(n6300), .Z(N101) );
  CEOX1 U9323 ( .A(N100), .B(mem_data1[82]), .Z(N8197) );
  CNR2X1 U9324 ( .A(n3838), .B(n6287), .Z(N100) );
  CEOX1 U9325 ( .A(N99), .B(mem_data1[81]), .Z(N8198) );
  CNR2X1 U9326 ( .A(n3840), .B(n6266), .Z(N99) );
  CEOX1 U9327 ( .A(N98), .B(mem_data1[80]), .Z(N8199) );
  CNR2X1 U9328 ( .A(n3842), .B(n6245), .Z(N98) );
  CEOX1 U9329 ( .A(N97), .B(mem_data1[79]), .Z(N8200) );
  CNR2X1 U9330 ( .A(n3837), .B(n6224), .Z(N97) );
  CEOX1 U9331 ( .A(N96), .B(mem_data1[78]), .Z(N8201) );
  CNR2X1 U9332 ( .A(n3847), .B(n6203), .Z(N96) );
  CEOX1 U9333 ( .A(N95), .B(mem_data1[77]), .Z(N8202) );
  CNR2X1 U9334 ( .A(n3841), .B(n6182), .Z(N95) );
  CEOX1 U9335 ( .A(N94), .B(mem_data1[76]), .Z(N8203) );
  CNR2X1 U9336 ( .A(n3851), .B(n6155), .Z(N94) );
  CEOX1 U9337 ( .A(N93), .B(mem_data1[75]), .Z(N8204) );
  CNR2X1 U9338 ( .A(n3849), .B(n6125), .Z(N93) );
  CEOX1 U9339 ( .A(N92), .B(mem_data1[74]), .Z(N8205) );
  CNR2X1 U9340 ( .A(n3852), .B(n6085), .Z(N92) );
  CEOX1 U9341 ( .A(N91), .B(mem_data1[73]), .Z(N8206) );
  CNR2X1 U9342 ( .A(n3851), .B(n6036), .Z(N91) );
  CEOX1 U9343 ( .A(N90), .B(mem_data1[72]), .Z(N8207) );
  CNR2X1 U9344 ( .A(n3849), .B(n6019), .Z(N90) );
  CEOX1 U9345 ( .A(N89), .B(mem_data1[71]), .Z(N8208) );
  CNR2X1 U9346 ( .A(n3849), .B(n6008), .Z(N89) );
  CEOX1 U9347 ( .A(N88), .B(mem_data1[70]), .Z(N8209) );
  CNR2X1 U9348 ( .A(n3848), .B(n5997), .Z(N88) );
  CEOX1 U9349 ( .A(N87), .B(mem_data1[69]), .Z(N8210) );
  CNR2X1 U9350 ( .A(n3847), .B(n5985), .Z(N87) );
  CEOX1 U9351 ( .A(N86), .B(mem_data1[68]), .Z(N8211) );
  CNR2X1 U9352 ( .A(n3846), .B(n5974), .Z(N86) );
  CEOX1 U9353 ( .A(N85), .B(mem_data1[67]), .Z(N8212) );
  CNR2X1 U9354 ( .A(n3845), .B(n5963), .Z(N85) );
  CEOX1 U9355 ( .A(N84), .B(mem_data1[66]), .Z(N8213) );
  CNR2X1 U9356 ( .A(n3844), .B(n5952), .Z(N84) );
  CEOX1 U9357 ( .A(N83), .B(mem_data1[65]), .Z(N8214) );
  CNR2X1 U9358 ( .A(n3843), .B(n5941), .Z(N83) );
  CEOX1 U9359 ( .A(N76), .B(mem_data1[58]), .Z(N8221) );
  CNR2X1 U9360 ( .A(n3844), .B(n5832), .Z(N76) );
  CEOX1 U9361 ( .A(N75), .B(mem_data1[57]), .Z(N8222) );
  CNR2X1 U9362 ( .A(n3838), .B(n5821), .Z(N75) );
  CEOX1 U9363 ( .A(N74), .B(mem_data1[56]), .Z(N8223) );
  CNR2X1 U9364 ( .A(n3848), .B(n5804), .Z(N74) );
  CEOX1 U9365 ( .A(N73), .B(mem_data1[55]), .Z(N8224) );
  CNR2X1 U9366 ( .A(n3842), .B(n5783), .Z(N73) );
  CEOX1 U9367 ( .A(N72), .B(mem_data1[54]), .Z(N8225) );
  CNR2X1 U9368 ( .A(n3845), .B(n5762), .Z(N72) );
  CEOX1 U9369 ( .A(N71), .B(mem_data1[53]), .Z(N8226) );
  CNR2X1 U9370 ( .A(n3846), .B(n5742), .Z(N71) );
  CEOX1 U9371 ( .A(N70), .B(mem_data1[52]), .Z(N8227) );
  CNR2X1 U9372 ( .A(n3836), .B(n5721), .Z(N70) );
  CEOX1 U9373 ( .A(N69), .B(mem_data1[51]), .Z(N8228) );
  CNR2X1 U9374 ( .A(n3850), .B(n5692), .Z(N69) );
  CEOX1 U9375 ( .A(N68), .B(mem_data1[50]), .Z(N8229) );
  CNR2X1 U9376 ( .A(n3853), .B(n5639), .Z(N68) );
  CEOX1 U9377 ( .A(N67), .B(mem_data1[49]), .Z(N8230) );
  CNR2X1 U9378 ( .A(n3843), .B(n5567), .Z(N67) );
  CEOX1 U9379 ( .A(N66), .B(mem_data1[48]), .Z(N8231) );
  CEOX1 U9380 ( .A(N65), .B(mem_data1[47]), .Z(N8232) );
  CNR2X1 U9381 ( .A(n3844), .B(n5462), .Z(N65) );
  CEOX1 U9382 ( .A(N63), .B(mem_data1[45]), .Z(N8234) );
  CNR2X1 U9383 ( .A(n3842), .B(n5440), .Z(N63) );
  CEOX1 U9384 ( .A(N62), .B(mem_data1[44]), .Z(N8235) );
  CNR2X1 U9385 ( .A(n3841), .B(n5429), .Z(N62) );
  CEOX1 U9386 ( .A(N61), .B(mem_data1[43]), .Z(N8236) );
  CNR2X1 U9387 ( .A(n3840), .B(n5418), .Z(N61) );
  CEOX1 U9388 ( .A(N60), .B(mem_data1[42]), .Z(N8237) );
  CNR2X1 U9389 ( .A(n3839), .B(n5407), .Z(N60) );
  CEOX1 U9390 ( .A(N59), .B(mem_data1[41]), .Z(N8238) );
  CNR2X1 U9391 ( .A(n3838), .B(n5396), .Z(N59) );
  CEOX1 U9392 ( .A(N58), .B(mem_data1[40]), .Z(N8239) );
  CNR2X1 U9393 ( .A(n3837), .B(n5385), .Z(N58) );
  CEOX1 U9394 ( .A(N57), .B(mem_data1[39]), .Z(N8240) );
  CNR2X1 U9395 ( .A(n3836), .B(n5373), .Z(N57) );
  CEOX1 U9396 ( .A(N56), .B(mem_data1[38]), .Z(N8241) );
  CNR2X1 U9397 ( .A(n3839), .B(n5362), .Z(N56) );
  CEOX1 U9398 ( .A(N55), .B(mem_data1[37]), .Z(N8242) );
  CNR2X1 U9399 ( .A(n3835), .B(n5347), .Z(N55) );
  CEOX1 U9400 ( .A(N51), .B(mem_data1[33]), .Z(N8246) );
  CNR2X1 U9401 ( .A(n3843), .B(n5276), .Z(N51) );
  CEOX1 U9402 ( .A(N50), .B(mem_data1[32]), .Z(N8247) );
  CNR2X1 U9403 ( .A(n3841), .B(n5265), .Z(N50) );
  CEOX1 U9404 ( .A(N49), .B(mem_data1[31]), .Z(N8248) );
  CNR2X1 U9405 ( .A(n3837), .B(n5254), .Z(N49) );
  CEOX1 U9406 ( .A(N48), .B(mem_data1[30]), .Z(N8249) );
  CNR2X1 U9407 ( .A(n3842), .B(n5233), .Z(N48) );
  CEOX1 U9408 ( .A(N47), .B(mem_data1[29]), .Z(N8250) );
  CNR2X1 U9409 ( .A(n3852), .B(n5211), .Z(N47) );
  CEOX1 U9410 ( .A(N46), .B(mem_data1[28]), .Z(N8251) );
  CNR2X1 U9411 ( .A(n3846), .B(n5190), .Z(N46) );
  CEOX1 U9412 ( .A(N45), .B(mem_data1[27]), .Z(N8252) );
  CNR2X1 U9413 ( .A(n3836), .B(n5170), .Z(N45) );
  CEOX1 U9414 ( .A(N44), .B(mem_data1[26]), .Z(N8253) );
  CNR2X1 U9415 ( .A(n3850), .B(n5147), .Z(N44) );
  CEOX1 U9416 ( .A(N43), .B(mem_data1[25]), .Z(N8254) );
  CNR2X1 U9417 ( .A(n3837), .B(n5112), .Z(N43) );
  CEOX1 U9418 ( .A(N42), .B(mem_data1[24]), .Z(N8255) );
  CNR2X1 U9419 ( .A(n3840), .B(n5047), .Z(N42) );
  CEOX1 U9420 ( .A(N41), .B(mem_data1[23]), .Z(N8256) );
  CNR2X1 U9421 ( .A(n3839), .B(n4977), .Z(N41) );
  CEOX1 U9422 ( .A(N40), .B(mem_data1[22]), .Z(N8257) );
  CNR2X1 U9423 ( .A(n3838), .B(n4922), .Z(N40) );
  CEOX1 U9424 ( .A(N39), .B(mem_data1[21]), .Z(N8258) );
  CNR2X1 U9425 ( .A(n3837), .B(n4903), .Z(N39) );
  CEOX1 U9426 ( .A(N38), .B(mem_data1[20]), .Z(N8259) );
  CNR2X1 U9427 ( .A(n3836), .B(n4892), .Z(N38) );
  CEOX1 U9428 ( .A(N37), .B(mem_data1[19]), .Z(N8260) );
  CNR2X1 U9429 ( .A(n3835), .B(n4880), .Z(N37) );
  CEOX1 U9430 ( .A(N36), .B(mem_data1[18]), .Z(N8261) );
  CNR2X1 U9431 ( .A(n3834), .B(n4867), .Z(N36) );
  CEOX1 U9432 ( .A(N35), .B(mem_data1[17]), .Z(N8262) );
  CNR2X1 U9433 ( .A(n3853), .B(n4846), .Z(N35) );
  CEOX1 U9434 ( .A(N34), .B(mem_data1[16]), .Z(N8263) );
  CNR2X1 U9435 ( .A(n3852), .B(n4825), .Z(N34) );
  CEOX1 U9436 ( .A(N33), .B(mem_data1[15]), .Z(N8264) );
  CNR2X1 U9437 ( .A(n3853), .B(n4805), .Z(N33) );
  CEOX1 U9438 ( .A(N694), .B(mem_data1[676]), .Z(N7603) );
  CNR2X1 U9439 ( .A(n3832), .B(n5959), .Z(N694) );
  CEOX1 U9440 ( .A(N1039), .B(mem_data1[1021]), .Z(N7258) );
  CNR2X1 U9441 ( .A(n3821), .B(n6388), .Z(N1039) );
  CEOX1 U9442 ( .A(N1038), .B(mem_data1[1020]), .Z(N7259) );
  CNR2X1 U9443 ( .A(n3818), .B(n6386), .Z(N1038) );
  CEOX1 U9444 ( .A(N1037), .B(mem_data1[1019]), .Z(N7260) );
  CNR2X1 U9445 ( .A(n3819), .B(n6384), .Z(N1037) );
  CEOX1 U9446 ( .A(N1036), .B(mem_data1[1018]), .Z(N7261) );
  CNR2X1 U9447 ( .A(n3820), .B(n6382), .Z(N1036) );
  CEOX1 U9448 ( .A(N1035), .B(mem_data1[1017]), .Z(N7262) );
  CNR2X1 U9449 ( .A(n3822), .B(n6379), .Z(N1035) );
  CEOX1 U9450 ( .A(N1034), .B(mem_data1[1016]), .Z(N7263) );
  CNR2X1 U9451 ( .A(n3823), .B(n6377), .Z(N1034) );
  CEOX1 U9452 ( .A(N1033), .B(mem_data1[1015]), .Z(N7264) );
  CNR2X1 U9453 ( .A(n3824), .B(n6375), .Z(N1033) );
  CEOX1 U9454 ( .A(N1032), .B(mem_data1[1014]), .Z(N7265) );
  CNR2X1 U9455 ( .A(n3825), .B(n6373), .Z(N1032) );
  CEOX1 U9456 ( .A(N1025), .B(mem_data1[1007]), .Z(N7272) );
  CNR2X1 U9457 ( .A(n3821), .B(n6358), .Z(N1025) );
  CEOX1 U9458 ( .A(N1024), .B(mem_data1[1006]), .Z(N7273) );
  CNR2X1 U9459 ( .A(n3822), .B(n6356), .Z(N1024) );
  CEOX1 U9460 ( .A(N1022), .B(mem_data1[1004]), .Z(N7275) );
  CNR2X1 U9461 ( .A(n3818), .B(n6352), .Z(N1022) );
  CEOX1 U9462 ( .A(N1019), .B(mem_data1[1001]), .Z(N7278) );
  CNR2X1 U9463 ( .A(n3816), .B(n6346), .Z(N1019) );
  CEOX1 U9464 ( .A(N1018), .B(mem_data1[1000]), .Z(N7279) );
  CNR2X1 U9465 ( .A(n3818), .B(n6344), .Z(N1018) );
  CEOX1 U9466 ( .A(N1017), .B(mem_data1[999]), .Z(N7280) );
  CNR2X1 U9467 ( .A(n3819), .B(n6511), .Z(N1017) );
  CEOX1 U9468 ( .A(N1015), .B(mem_data1[997]), .Z(N7282) );
  CNR2X1 U9469 ( .A(n3823), .B(n6509), .Z(N1015) );
  CEOX1 U9470 ( .A(N1014), .B(mem_data1[996]), .Z(N7283) );
  CNR2X1 U9471 ( .A(n3822), .B(n6508), .Z(N1014) );
  CEOX1 U9472 ( .A(N1013), .B(mem_data1[995]), .Z(N7284) );
  CNR2X1 U9473 ( .A(n3827), .B(n6507), .Z(N1013) );
  CEOX1 U9474 ( .A(N1012), .B(mem_data1[994]), .Z(N7285) );
  CNR2X1 U9475 ( .A(n3826), .B(n6506), .Z(N1012) );
  CEOX1 U9476 ( .A(N1011), .B(mem_data1[993]), .Z(N7286) );
  CNR2X1 U9477 ( .A(n3825), .B(n6505), .Z(N1011) );
  CEOX1 U9478 ( .A(N1010), .B(mem_data1[992]), .Z(N7287) );
  CNR2X1 U9479 ( .A(n3830), .B(n6504), .Z(N1010) );
  CEOX1 U9480 ( .A(N978), .B(mem_data1[960]), .Z(N7319) );
  CNR2X1 U9481 ( .A(n3824), .B(n6465), .Z(N978) );
  CEOX1 U9482 ( .A(N946), .B(mem_data1[928]), .Z(N7351) );
  CNR2X1 U9483 ( .A(n3817), .B(n6429), .Z(N946) );
  CEOX1 U9484 ( .A(N914), .B(mem_data1[896]), .Z(N7383) );
  CNR2X1 U9485 ( .A(n3818), .B(n6393), .Z(N914) );
  CEOX1 U9486 ( .A(N882), .B(mem_data1[864]), .Z(N7415) );
  CNR2X1 U9487 ( .A(n3844), .B(n6504), .Z(N882) );
  CEOX1 U9488 ( .A(N850), .B(mem_data1[832]), .Z(N7447) );
  CNR2X1 U9489 ( .A(n3841), .B(n6465), .Z(N850) );
  CEOX1 U9490 ( .A(N818), .B(mem_data1[800]), .Z(N7479) );
  CNR2X1 U9491 ( .A(n3851), .B(n6429), .Z(N818) );
  CEOX1 U9492 ( .A(N786), .B(mem_data1[768]), .Z(N7511) );
  CNR2X1 U9493 ( .A(n3853), .B(n6393), .Z(N786) );
  CEOX1 U9494 ( .A(N771), .B(mem_data1[753]), .Z(N7526) );
  CEOX1 U9495 ( .A(N770), .B(mem_data1[752]), .Z(N7527) );
  CEOX1 U9496 ( .A(N760), .B(mem_data1[742]), .Z(N7537) );
  CEOX1 U9497 ( .A(N754), .B(mem_data1[736]), .Z(N7543) );
  CNR2X1 U9498 ( .A(n3826), .B(n6026), .Z(N754) );
  CEOX1 U9499 ( .A(N748), .B(mem_data1[730]), .Z(N7549) );
  CNR2X1 U9500 ( .A(n3816), .B(n6020), .Z(N748) );
  CEOX1 U9501 ( .A(N738), .B(mem_data1[720]), .Z(N7559) );
  CNR2X1 U9502 ( .A(n3825), .B(n6009), .Z(N738) );
  CEOX1 U9503 ( .A(N734), .B(mem_data1[716]), .Z(N7563) );
  CNR2X1 U9504 ( .A(n3821), .B(n6004), .Z(N734) );
  CEOX1 U9505 ( .A(N733), .B(mem_data1[715]), .Z(N7564) );
  CNR2X1 U9506 ( .A(n3817), .B(n6003), .Z(N733) );
  CEOX1 U9507 ( .A(N702), .B(mem_data1[684]), .Z(N7595) );
  CNR2X1 U9508 ( .A(n3817), .B(n5968), .Z(N702) );
  CEOX1 U9509 ( .A(N700), .B(mem_data1[682]), .Z(N7597) );
  CNR2X1 U9510 ( .A(n3827), .B(n5966), .Z(N700) );
  CEOX1 U9511 ( .A(N696), .B(mem_data1[678]), .Z(N7601) );
  CNR2X1 U9512 ( .A(n3815), .B(n5961), .Z(N696) );
  CEOX1 U9513 ( .A(N690), .B(mem_data1[672]), .Z(N7607) );
  CNR2X1 U9514 ( .A(n3830), .B(n5955), .Z(N690) );
  CEOX1 U9515 ( .A(N684), .B(mem_data1[666]), .Z(N7613) );
  CNR2X1 U9516 ( .A(n3831), .B(n5948), .Z(N684) );
  CEOX1 U9517 ( .A(N674), .B(mem_data1[656]), .Z(N7623) );
  CNR2X1 U9518 ( .A(n3828), .B(n5937), .Z(N674) );
  CEOX1 U9519 ( .A(N669), .B(mem_data1[651]), .Z(N7628) );
  CNR2X1 U9520 ( .A(n3821), .B(n5932), .Z(N669) );
  CEOX1 U9521 ( .A(N662), .B(mem_data1[644]), .Z(N7635) );
  CNR2X1 U9522 ( .A(n3816), .B(n5924), .Z(N662) );
  CEOX1 U9523 ( .A(N632), .B(mem_data1[614]), .Z(N7665) );
  CEOX1 U9524 ( .A(N626), .B(mem_data1[608]), .Z(N7671) );
  CNR2X1 U9525 ( .A(n3838), .B(n6026), .Z(N626) );
  CEOX1 U9526 ( .A(N623), .B(mem_data1[605]), .Z(N7674) );
  CNR2X1 U9527 ( .A(n3850), .B(n6023), .Z(N623) );
  CEOX1 U9528 ( .A(N620), .B(mem_data1[602]), .Z(N7677) );
  CNR2X1 U9529 ( .A(n3848), .B(n6020), .Z(N620) );
  CEOX1 U9530 ( .A(N610), .B(mem_data1[592]), .Z(N7687) );
  CNR2X1 U9531 ( .A(n3846), .B(n6009), .Z(N610) );
  CEOX1 U9532 ( .A(N606), .B(mem_data1[588]), .Z(N7691) );
  CNR2X1 U9533 ( .A(n3842), .B(n6004), .Z(N606) );
  CEOX1 U9534 ( .A(N605), .B(mem_data1[587]), .Z(N7692) );
  CNR2X1 U9535 ( .A(n3847), .B(n6003), .Z(N605) );
  CEOX1 U9536 ( .A(N594), .B(mem_data1[576]), .Z(N7703) );
  CNR2X1 U9537 ( .A(n3834), .B(n5991), .Z(N594) );
  CEOX1 U9538 ( .A(N574), .B(mem_data1[556]), .Z(N7723) );
  CNR2X1 U9539 ( .A(n3838), .B(n5968), .Z(N574) );
  CEOX1 U9540 ( .A(N572), .B(mem_data1[554]), .Z(N7725) );
  CNR2X1 U9541 ( .A(n3837), .B(n5966), .Z(N572) );
  CEOX1 U9542 ( .A(N568), .B(mem_data1[550]), .Z(N7729) );
  CNR2X1 U9543 ( .A(n3841), .B(n5961), .Z(N568) );
  CEOX1 U9544 ( .A(N562), .B(mem_data1[544]), .Z(N7735) );
  CNR2X1 U9545 ( .A(n3851), .B(n5955), .Z(N562) );
  CEOX1 U9546 ( .A(N556), .B(mem_data1[538]), .Z(N7741) );
  CNR2X1 U9547 ( .A(n3844), .B(n5948), .Z(N556) );
  CEOX1 U9548 ( .A(N546), .B(mem_data1[528]), .Z(N7751) );
  CNR2X1 U9549 ( .A(n3839), .B(n5937), .Z(N546) );
  CEOX1 U9550 ( .A(N541), .B(mem_data1[523]), .Z(N7756) );
  CNR2X1 U9551 ( .A(n3834), .B(n5932), .Z(N541) );
  CEOX1 U9552 ( .A(N534), .B(mem_data1[516]), .Z(N7763) );
  CNR2X1 U9553 ( .A(n3847), .B(n5924), .Z(N534) );
  CEOX1 U9554 ( .A(N530), .B(mem_data1[512]), .Z(N7767) );
  CNR2X1 U9555 ( .A(n3834), .B(n5920), .Z(N530) );
  CEOX1 U9556 ( .A(N1040), .B(mem_data1[1022]), .Z(N7257) );
  CNR2X1 U9557 ( .A(n3816), .B(n6390), .Z(N1040) );
  CNR2X1 U9558 ( .A(n4434), .B(reqin0), .Z(n79) );
  CEOX1 U9559 ( .A(N1041), .B(mem_data1[1023]), .Z(N7256) );
  CNR2X1 U9560 ( .A(n3817), .B(n6392), .Z(N1041) );
  CEOX1 U9561 ( .A(N399), .B(mem_data1[381]), .Z(N7898) );
  CEOX1 U9562 ( .A(N375), .B(mem_data1[357]), .Z(N7922) );
  CEOX1 U9563 ( .A(N505), .B(mem_data1[487]), .Z(N7792) );
  CEOX1 U9564 ( .A(N503), .B(mem_data1[485]), .Z(N7794) );
  CEOX1 U9565 ( .A(N401), .B(mem_data1[383]), .Z(N7896) );
  CEOX1 U9566 ( .A(N273), .B(mem_data1[255]), .Z(N8024) );
  CEOX1 U9567 ( .A(N271), .B(mem_data1[253]), .Z(N8026) );
  CEOX1 U9568 ( .A(N518), .B(mem_data1[500]), .Z(N7779) );
  CEOX1 U9569 ( .A(N515), .B(mem_data1[497]), .Z(N7782) );
  CEOX1 U9570 ( .A(N496), .B(mem_data1[478]), .Z(N7801) );
  CNR2X1 U9571 ( .A(n3823), .B(n5460), .Z(N496) );
  CEOX1 U9572 ( .A(N484), .B(mem_data1[466]), .Z(N7813) );
  CNR2X1 U9573 ( .A(n3824), .B(n5447), .Z(N484) );
  CEOX1 U9574 ( .A(N474), .B(mem_data1[456]), .Z(N7823) );
  CNR2X1 U9575 ( .A(n3829), .B(n5436), .Z(N474) );
  CEOX1 U9576 ( .A(N422), .B(mem_data1[404]), .Z(N7875) );
  CNR2X1 U9577 ( .A(n3831), .B(n5379), .Z(N422) );
  CEOX1 U9578 ( .A(N414), .B(mem_data1[396]), .Z(N7883) );
  CNR2X1 U9579 ( .A(n3821), .B(n5369), .Z(N414) );
  CEOX1 U9580 ( .A(N410), .B(mem_data1[392]), .Z(N7887) );
  CNR2X1 U9581 ( .A(n3817), .B(n5365), .Z(N410) );
  CEOX1 U9582 ( .A(N402), .B(mem_data1[384]), .Z(N7895) );
  CNR2X1 U9583 ( .A(n3830), .B(n5356), .Z(N402) );
  CEOX1 U9584 ( .A(N368), .B(mem_data1[350]), .Z(N7929) );
  CNR2X1 U9585 ( .A(n3842), .B(n5460), .Z(N368) );
  CEOX1 U9586 ( .A(N358), .B(mem_data1[340]), .Z(N7939) );
  CNR2X1 U9587 ( .A(n3844), .B(n5449), .Z(N358) );
  CEOX1 U9588 ( .A(N354), .B(mem_data1[336]), .Z(N7943) );
  CNR2X1 U9589 ( .A(n3840), .B(n5445), .Z(N354) );
  CEOX1 U9590 ( .A(N350), .B(mem_data1[332]), .Z(N7947) );
  CNR2X1 U9591 ( .A(n3841), .B(n5441), .Z(N350) );
  CEOX1 U9592 ( .A(N346), .B(mem_data1[328]), .Z(N7951) );
  CNR2X1 U9593 ( .A(n3836), .B(n5436), .Z(N346) );
  CEOX1 U9594 ( .A(N338), .B(mem_data1[320]), .Z(N7959) );
  CNR2X1 U9595 ( .A(n3848), .B(n5427), .Z(N338) );
  CEOX1 U9596 ( .A(N304), .B(mem_data1[286]), .Z(N7993) );
  CNR2X1 U9597 ( .A(n3842), .B(n5390), .Z(N304) );
  CEOX1 U9598 ( .A(N294), .B(mem_data1[276]), .Z(N8003) );
  CNR2X1 U9599 ( .A(n3838), .B(n5379), .Z(N294) );
  CEOX1 U9600 ( .A(N290), .B(mem_data1[272]), .Z(N8007) );
  CNR2X1 U9601 ( .A(n3853), .B(n5375), .Z(N290) );
  CEOX1 U9602 ( .A(N286), .B(mem_data1[268]), .Z(N8011) );
  CNR2X1 U9603 ( .A(n3848), .B(n5369), .Z(N286) );
  CEOX1 U9604 ( .A(N282), .B(mem_data1[264]), .Z(N8015) );
  CNR2X1 U9605 ( .A(n3845), .B(n5365), .Z(N282) );
  CEOX1 U9606 ( .A(N274), .B(mem_data1[256]), .Z(N8023) );
  CNR2X1 U9607 ( .A(n3841), .B(n5356), .Z(N274) );
  CEOX1 U9608 ( .A(N251), .B(mem_data1[233]), .Z(N8046) );
  CEOX1 U9609 ( .A(N182), .B(mem_data1[164]), .Z(N8115) );
  CEOX1 U9610 ( .A(N146), .B(mem_data1[128]), .Z(N8151) );
  CNR2X1 U9611 ( .A(n3827), .B(n4738), .Z(N146) );
  CEOX1 U9612 ( .A(N129), .B(mem_data1[111]), .Z(N8168) );
  CEOX1 U9613 ( .A(N123), .B(mem_data1[105]), .Z(N8174) );
  CEOX1 U9614 ( .A(N113), .B(mem_data1[95]), .Z(N8184) );
  CNR2X1 U9615 ( .A(n3851), .B(n6464), .Z(N113) );
  CEOX1 U9616 ( .A(N82), .B(mem_data1[64]), .Z(N8215) );
  CNR2X1 U9617 ( .A(n3842), .B(n5930), .Z(N82) );
  CEOX1 U9618 ( .A(N54), .B(mem_data1[36]), .Z(N8243) );
  CEOX1 U9619 ( .A(N370), .B(mem_data1[352]), .Z(N7927) );
  CNR2X1 U9620 ( .A(n3852), .B(n5463), .Z(N370) );
  CEOX1 U9621 ( .A(N516), .B(mem_data1[498]), .Z(N7781) );
  CEOX1 U9622 ( .A(N498), .B(mem_data1[480]), .Z(N7799) );
  CNR2X1 U9623 ( .A(n3819), .B(n5463), .Z(N498) );
  CEOX1 U9624 ( .A(N494), .B(mem_data1[476]), .Z(N7803) );
  CNR2X1 U9625 ( .A(n3832), .B(n5458), .Z(N494) );
  CEOX1 U9626 ( .A(N480), .B(mem_data1[462]), .Z(N7817) );
  CNR2X1 U9627 ( .A(n3818), .B(n5443), .Z(N480) );
  CEOX1 U9628 ( .A(N470), .B(mem_data1[452]), .Z(N7827) );
  CNR2X1 U9629 ( .A(n3827), .B(n5432), .Z(N470) );
  CEOX1 U9630 ( .A(N430), .B(mem_data1[412]), .Z(N7867) );
  CNR2X1 U9631 ( .A(n3815), .B(n5388), .Z(N430) );
  CEOX1 U9632 ( .A(N416), .B(mem_data1[398]), .Z(N7881) );
  CNR2X1 U9633 ( .A(n3825), .B(n5371), .Z(N416) );
  CEOX1 U9634 ( .A(N412), .B(mem_data1[394]), .Z(N7885) );
  CNR2X1 U9635 ( .A(n3818), .B(n5367), .Z(N412) );
  CEOX1 U9636 ( .A(N408), .B(mem_data1[390]), .Z(N7889) );
  CNR2X1 U9637 ( .A(n3831), .B(n5363), .Z(N408) );
  CEOX1 U9638 ( .A(N366), .B(mem_data1[348]), .Z(N7931) );
  CNR2X1 U9639 ( .A(n3842), .B(n5458), .Z(N366) );
  CEOX1 U9640 ( .A(N356), .B(mem_data1[338]), .Z(N7941) );
  CNR2X1 U9641 ( .A(n3838), .B(n5447), .Z(N356) );
  CEOX1 U9642 ( .A(N352), .B(mem_data1[334]), .Z(N7945) );
  CNR2X1 U9643 ( .A(n3838), .B(n5443), .Z(N352) );
  CEOX1 U9644 ( .A(N348), .B(mem_data1[330]), .Z(N7949) );
  CNR2X1 U9645 ( .A(n3847), .B(n5438), .Z(N348) );
  CEOX1 U9646 ( .A(N342), .B(mem_data1[324]), .Z(N7955) );
  CNR2X1 U9647 ( .A(n3852), .B(n5432), .Z(N342) );
  CEOX1 U9648 ( .A(N329), .B(mem_data1[311]), .Z(N7968) );
  CNR2X1 U9649 ( .A(n3840), .B(n5417), .Z(N329) );
  CEOX1 U9650 ( .A(N306), .B(mem_data1[288]), .Z(N7991) );
  CNR2X1 U9651 ( .A(n3844), .B(n5392), .Z(N306) );
  CEOX1 U9652 ( .A(N302), .B(mem_data1[284]), .Z(N7995) );
  CNR2X1 U9653 ( .A(n3840), .B(n5388), .Z(N302) );
  CEOX1 U9654 ( .A(N292), .B(mem_data1[274]), .Z(N8005) );
  CNR2X1 U9655 ( .A(n3835), .B(n5377), .Z(N292) );
  CEOX1 U9656 ( .A(N284), .B(mem_data1[266]), .Z(N8013) );
  CNR2X1 U9657 ( .A(n3846), .B(n5367), .Z(N284) );
  CEOX1 U9658 ( .A(N278), .B(mem_data1[260]), .Z(N8019) );
  CNR2X1 U9659 ( .A(n3837), .B(n5360), .Z(N278) );
  CEOX1 U9660 ( .A(N255), .B(mem_data1[237]), .Z(N8042) );
  CEOX1 U9661 ( .A(N244), .B(mem_data1[226]), .Z(N8053) );
  CEOX1 U9662 ( .A(N239), .B(mem_data1[221]), .Z(N8058) );
  CNR2X1 U9663 ( .A(n3826), .B(n6442), .Z(N239) );
  CEOX1 U9664 ( .A(N206), .B(mem_data1[188]), .Z(N8091) );
  CNR2X1 U9665 ( .A(n3831), .B(n5856), .Z(N206) );
  CEOX1 U9666 ( .A(N126), .B(mem_data1[108]), .Z(N8171) );
  CEOX1 U9667 ( .A(N114), .B(mem_data1[96]), .Z(N8183) );
  CNR2X1 U9668 ( .A(n3852), .B(n6475), .Z(N114) );
  CEOX1 U9669 ( .A(N111), .B(mem_data1[93]), .Z(N8186) );
  CNR2X1 U9670 ( .A(n3849), .B(n6442), .Z(N111) );
  CEOX1 U9671 ( .A(N77), .B(mem_data1[59]), .Z(N8220) );
  CNR2X1 U9672 ( .A(n3834), .B(n5843), .Z(N77) );
  CEOX1 U9673 ( .A(N52), .B(mem_data1[34]), .Z(N8245) );
  CNR2X1 U9674 ( .A(n3851), .B(n5287), .Z(N52) );
  CEOX1 U9675 ( .A(N32), .B(mem_data1[14]), .Z(N8265) );
  CNR2X1 U9676 ( .A(n3853), .B(n4784), .Z(N32) );
  CEOX1 U9677 ( .A(N434), .B(mem_data1[416]), .Z(N7863) );
  CNR2X1 U9678 ( .A(n3822), .B(n5392), .Z(N434) );
  CEOX1 U9679 ( .A(N450), .B(mem_data1[432]), .Z(N7847) );
  CNR2X1 U9680 ( .A(n3831), .B(n5410), .Z(N450) );
  CEOX1 U9681 ( .A(N482), .B(mem_data1[464]), .Z(N7815) );
  CNR2X1 U9682 ( .A(n3820), .B(n5445), .Z(N482) );
  CEOX1 U9683 ( .A(N472), .B(mem_data1[454]), .Z(N7825) );
  CNR2X1 U9684 ( .A(n3831), .B(n5434), .Z(N472) );
  CNR2X1 U9685 ( .A(n3815), .B(n5412), .Z(N452) );
  CEOX1 U9686 ( .A(N447), .B(mem_data1[429]), .Z(N7850) );
  CNR2X1 U9687 ( .A(n3828), .B(n5406), .Z(N447) );
  CEOX1 U9688 ( .A(N432), .B(mem_data1[414]), .Z(N7865) );
  CNR2X1 U9689 ( .A(n3825), .B(n5390), .Z(N432) );
  CEOX1 U9690 ( .A(N420), .B(mem_data1[402]), .Z(N7877) );
  CNR2X1 U9691 ( .A(n3827), .B(n5377), .Z(N420) );
  CEOX1 U9692 ( .A(N388), .B(mem_data1[370]), .Z(N7909) );
  CEOX1 U9693 ( .A(N386), .B(mem_data1[368]), .Z(N7911) );
  CEOX1 U9694 ( .A(N344), .B(mem_data1[326]), .Z(N7953) );
  CNR2X1 U9695 ( .A(n3834), .B(n5434), .Z(N344) );
  CEOX1 U9696 ( .A(N322), .B(mem_data1[304]), .Z(N7975) );
  CNR2X1 U9697 ( .A(n3836), .B(n5410), .Z(N322) );
  CEOX1 U9698 ( .A(N319), .B(mem_data1[301]), .Z(N7978) );
  CNR2X1 U9699 ( .A(n3836), .B(n5406), .Z(N319) );
  CEOX1 U9700 ( .A(N280), .B(mem_data1[262]), .Z(N8017) );
  CNR2X1 U9701 ( .A(n3843), .B(n5363), .Z(N280) );
  CEOX1 U9702 ( .A(N260), .B(mem_data1[242]), .Z(N8037) );
  CEOX1 U9703 ( .A(N258), .B(mem_data1[240]), .Z(N8039) );
  CEOX1 U9704 ( .A(N246), .B(mem_data1[228]), .Z(N8051) );
  CEOX1 U9705 ( .A(N142), .B(mem_data1[124]), .Z(N8155) );
  CEOX1 U9706 ( .A(N118), .B(mem_data1[100]), .Z(N8179) );
  CND2X1 U9707 ( .A(n4814), .B(n3723), .Z(n4518) );
  CEOX1 U9708 ( .A(N116), .B(mem_data1[98]), .Z(N8181) );
  CEOX1 U9709 ( .A(N80), .B(mem_data1[62]), .Z(N8217) );
  CNR2X1 U9710 ( .A(n3840), .B(n5898), .Z(N80) );
  CEOX1 U9711 ( .A(N369), .B(mem_data1[351]), .Z(N7928) );
  CNR2X1 U9712 ( .A(n3852), .B(n5461), .Z(N369) );
  CEOX1 U9713 ( .A(N497), .B(mem_data1[479]), .Z(N7800) );
  CNR2X1 U9714 ( .A(n3827), .B(n5461), .Z(N497) );
  CEOX1 U9715 ( .A(N305), .B(mem_data1[287]), .Z(N7992) );
  CNR2X1 U9716 ( .A(n3843), .B(n5391), .Z(N305) );
  CEOX1 U9717 ( .A(N192), .B(mem_data1[174]), .Z(N8105) );
  CNR2X1 U9718 ( .A(n3820), .B(n5451), .Z(N192) );
  CEOX1 U9719 ( .A(N64), .B(mem_data1[46]), .Z(N8233) );
  CNR2X1 U9720 ( .A(n3843), .B(n5451), .Z(N64) );
  CEOX1 U9721 ( .A(N328), .B(mem_data1[310]), .Z(N7969) );
  CNR2X1 U9722 ( .A(n3843), .B(n5416), .Z(N328) );
  CEOX1 U9723 ( .A(N208), .B(mem_data1[190]), .Z(N8089) );
  CNR2X1 U9724 ( .A(n3815), .B(n5898), .Z(N208) );
  CEOX1 U9725 ( .A(N289), .B(mem_data1[271]), .Z(N8008) );
  CNR2X1 U9726 ( .A(n3852), .B(n5372), .Z(N289) );
  CEOX1 U9727 ( .A(N180), .B(mem_data1[162]), .Z(N8117) );
  CNR2X1 U9728 ( .A(n3823), .B(n5287), .Z(N180) );
  CEOX1 U9729 ( .A(mem_data1[445]), .B(N463), .Z(N7834) );
  CNR2IX1 U9730 ( .B(n3839), .A(n5424), .Z(N463) );
  CEOX1 U9731 ( .A(mem_data1[447]), .B(N465), .Z(N7832) );
  CNR2IX1 U9732 ( .B(n3840), .A(n5426), .Z(N465) );
  CEOX1 U9733 ( .A(N176), .B(mem_data1[158]), .Z(N8121) );
  CNR2X1 U9734 ( .A(n3832), .B(n5233), .Z(N176) );
  CEOX1 U9735 ( .A(mem_data1[296]), .B(N314), .Z(N7983) );
  CNR2IX1 U9736 ( .B(n3832), .A(n5401), .Z(N314) );
  CEOX1 U9737 ( .A(mem_data1[303]), .B(N321), .Z(N7976) );
  CNR2IX1 U9738 ( .B(n3827), .A(n5409), .Z(N321) );
  CEOX1 U9739 ( .A(mem_data1[305]), .B(N323), .Z(N7974) );
  CNR2IX1 U9740 ( .B(n3829), .A(n5411), .Z(N323) );
  CEOX1 U9741 ( .A(N457), .B(mem_data1[439]), .Z(N7840) );
  CNR2X1 U9742 ( .A(n3816), .B(n5417), .Z(N457) );
  CEOX1 U9743 ( .A(mem_data1[430]), .B(N448), .Z(N7849) );
  CNR2IX1 U9744 ( .B(n3845), .A(n5408), .Z(N448) );
  CEOX1 U9745 ( .A(mem_data1[427]), .B(N445), .Z(N7852) );
  CNR2IX1 U9746 ( .B(n3839), .A(n5404), .Z(N445) );
  CEOX1 U9747 ( .A(N442), .B(mem_data1[424]), .Z(N7855) );
  CNR2X1 U9748 ( .A(n3827), .B(n5401), .Z(N442) );
  CEOX1 U9749 ( .A(N181), .B(mem_data1[163]), .Z(N8116) );
  CNR2X1 U9750 ( .A(n3833), .B(n5305), .Z(N181) );
  CEOX1 U9751 ( .A(N53), .B(mem_data1[35]), .Z(N8244) );
  CNR2X1 U9752 ( .A(n3853), .B(n5305), .Z(N53) );
  CEOX1 U9753 ( .A(N240), .B(mem_data1[222]), .Z(N8057) );
  CNR2X1 U9754 ( .A(n3818), .B(n6453), .Z(N240) );
  CEOX1 U9755 ( .A(N137), .B(mem_data1[119]), .Z(N8160) );
  CEOX1 U9756 ( .A(N396), .B(mem_data1[378]), .Z(N7901) );
  CEOX1 U9757 ( .A(N317), .B(mem_data1[299]), .Z(N7980) );
  CNR2IX1 U9758 ( .B(n3830), .A(n5404), .Z(N317) );
  CEOX1 U9759 ( .A(N141), .B(mem_data1[123]), .Z(N8156) );
  CEOX1 U9760 ( .A(N139), .B(mem_data1[121]), .Z(N8158) );
  CEOX1 U9761 ( .A(N310), .B(mem_data1[292]), .Z(N7987) );
  CNR2X1 U9762 ( .A(n3849), .B(n5397), .Z(N310) );
  CEOX1 U9763 ( .A(mem_data1[294]), .B(N312), .Z(N7985) );
  CNR2IX1 U9764 ( .B(n3819), .A(n5399), .Z(N312) );
  CEOX1 U9765 ( .A(mem_data1[290]), .B(N308), .Z(N7989) );
  CNR2IX1 U9766 ( .B(n3820), .A(n5394), .Z(N308) );
  CEOX1 U9767 ( .A(N333), .B(mem_data1[315]), .Z(N7964) );
  CNR2X1 U9768 ( .A(n3846), .B(n5422), .Z(N333) );
  CEOX1 U9769 ( .A(mem_data1[317]), .B(N335), .Z(N7962) );
  CNR2IX1 U9770 ( .B(n3815), .A(n5424), .Z(N335) );
  CEOX1 U9771 ( .A(N512), .B(mem_data1[494]), .Z(N7785) );
  CEOX1 U9772 ( .A(N495), .B(mem_data1[477]), .Z(N7802) );
  CNR2IX1 U9773 ( .B(n3839), .A(n5459), .Z(N495) );
  CEOX1 U9774 ( .A(N483), .B(mem_data1[465]), .Z(N7814) );
  CNR2X1 U9775 ( .A(n3819), .B(n5446), .Z(N483) );
  CEOX1 U9776 ( .A(N481), .B(mem_data1[463]), .Z(N7816) );
  CNR2X1 U9777 ( .A(n3821), .B(n5444), .Z(N481) );
  CEOX1 U9778 ( .A(N473), .B(mem_data1[455]), .Z(N7824) );
  CNR2X1 U9779 ( .A(n3830), .B(n5435), .Z(N473) );
  CEOX1 U9780 ( .A(N471), .B(mem_data1[453]), .Z(N7826) );
  CNR2X1 U9781 ( .A(n3826), .B(n5433), .Z(N471) );
  CEOX1 U9782 ( .A(N458), .B(mem_data1[440]), .Z(N7839) );
  CNR2IX1 U9783 ( .B(n3841), .A(n5419), .Z(N458) );
  CEOX1 U9784 ( .A(N456), .B(mem_data1[438]), .Z(N7841) );
  CNR2X1 U9785 ( .A(n3817), .B(n5416), .Z(N456) );
  CEOX1 U9786 ( .A(mem_data1[435]), .B(N453), .Z(N7844) );
  CNR2IX1 U9787 ( .B(n3845), .A(n5413), .Z(N453) );
  CEOX1 U9788 ( .A(mem_data1[433]), .B(N451), .Z(N7846) );
  CNR2IX1 U9789 ( .B(n3842), .A(n5411), .Z(N451) );
  CEOX1 U9790 ( .A(mem_data1[431]), .B(N449), .Z(N7848) );
  CNR2IX1 U9791 ( .B(n3842), .A(n5409), .Z(N449) );
  CEOX1 U9792 ( .A(N446), .B(mem_data1[428]), .Z(N7851) );
  CNR2X1 U9793 ( .A(n3829), .B(n5405), .Z(N446) );
  CEOX1 U9794 ( .A(N444), .B(mem_data1[426]), .Z(N7853) );
  CNR2X1 U9795 ( .A(n3829), .B(n5403), .Z(N444) );
  CEOX1 U9796 ( .A(N443), .B(mem_data1[425]), .Z(N7854) );
  CNR2X1 U9797 ( .A(n3826), .B(n5402), .Z(N443) );
  CEOX1 U9798 ( .A(mem_data1[423]), .B(N441), .Z(N7856) );
  CNR2IX1 U9799 ( .B(n3845), .A(n5400), .Z(N441) );
  CEOX1 U9800 ( .A(mem_data1[422]), .B(N440), .Z(N7857) );
  CNR2IX1 U9801 ( .B(n3840), .A(n5399), .Z(N440) );
  CEOX1 U9802 ( .A(mem_data1[421]), .B(N439), .Z(N7858) );
  CNR2IX1 U9803 ( .B(n3839), .A(n5398), .Z(N439) );
  CEOX1 U9804 ( .A(N438), .B(mem_data1[420]), .Z(N7859) );
  CNR2X1 U9805 ( .A(n3821), .B(n5397), .Z(N438) );
  CEOX1 U9806 ( .A(mem_data1[418]), .B(N436), .Z(N7861) );
  CNR2IX1 U9807 ( .B(n3845), .A(n5394), .Z(N436) );
  CEOX1 U9808 ( .A(N433), .B(mem_data1[415]), .Z(N7864) );
  CNR2X1 U9809 ( .A(n3824), .B(n5391), .Z(N433) );
  CEOX1 U9810 ( .A(N421), .B(mem_data1[403]), .Z(N7876) );
  CNR2X1 U9811 ( .A(n3826), .B(n5378), .Z(N421) );
  CEOX1 U9812 ( .A(N419), .B(mem_data1[401]), .Z(N7878) );
  CNR2X1 U9813 ( .A(n3828), .B(n5376), .Z(N419) );
  CEOX1 U9814 ( .A(N418), .B(mem_data1[400]), .Z(N7879) );
  CNR2X1 U9815 ( .A(n3823), .B(n5375), .Z(N418) );
  CEOX1 U9816 ( .A(N417), .B(mem_data1[399]), .Z(N7880) );
  CNR2X1 U9817 ( .A(n3824), .B(n5372), .Z(N417) );
  CEOX1 U9818 ( .A(N413), .B(mem_data1[395]), .Z(N7884) );
  CNR2X1 U9819 ( .A(n3822), .B(n5368), .Z(N413) );
  CEOX1 U9820 ( .A(N409), .B(mem_data1[391]), .Z(N7888) );
  CNR2X1 U9821 ( .A(n3820), .B(n5364), .Z(N409) );
  CEOX1 U9822 ( .A(N400), .B(mem_data1[382]), .Z(N7897) );
  CEOX1 U9823 ( .A(N383), .B(mem_data1[365]), .Z(N7914) );
  CEOX1 U9824 ( .A(N367), .B(mem_data1[349]), .Z(N7930) );
  CNR2X1 U9825 ( .A(n3850), .B(n5459), .Z(N367) );
  CEOX1 U9826 ( .A(N357), .B(mem_data1[339]), .Z(N7940) );
  CNR2X1 U9827 ( .A(n3842), .B(n5448), .Z(N357) );
  CEOX1 U9828 ( .A(N353), .B(mem_data1[335]), .Z(N7944) );
  CNR2X1 U9829 ( .A(n3839), .B(n5444), .Z(N353) );
  CEOX1 U9830 ( .A(N349), .B(mem_data1[331]), .Z(N7948) );
  CNR2X1 U9831 ( .A(n3848), .B(n5439), .Z(N349) );
  CEOX1 U9832 ( .A(N345), .B(mem_data1[327]), .Z(N7952) );
  CNR2X1 U9833 ( .A(n3835), .B(n5435), .Z(N345) );
  CEOX1 U9834 ( .A(N343), .B(mem_data1[325]), .Z(N7954) );
  CNR2X1 U9835 ( .A(n3853), .B(n5433), .Z(N343) );
  CEOX1 U9836 ( .A(mem_data1[319]), .B(N337), .Z(N7960) );
  CNR2IX1 U9837 ( .B(n3823), .A(n5426), .Z(N337) );
  CEOX1 U9838 ( .A(N336), .B(mem_data1[318]), .Z(N7961) );
  CNR2X1 U9839 ( .A(n3846), .B(n5425), .Z(N336) );
  CEOX1 U9840 ( .A(N334), .B(mem_data1[316]), .Z(N7963) );
  CNR2X1 U9841 ( .A(n3844), .B(n5423), .Z(N334) );
  CEOX1 U9842 ( .A(N332), .B(mem_data1[314]), .Z(N7965) );
  CNR2X1 U9843 ( .A(n3840), .B(n5421), .Z(N332) );
  CEOX1 U9844 ( .A(N331), .B(mem_data1[313]), .Z(N7966) );
  CNR2X1 U9845 ( .A(n3845), .B(n5420), .Z(N331) );
  CEOX1 U9846 ( .A(N330), .B(mem_data1[312]), .Z(N7967) );
  CNR2X1 U9847 ( .A(n3844), .B(n5419), .Z(N330) );
  CEOX1 U9848 ( .A(N327), .B(mem_data1[309]), .Z(N7970) );
  CNR2X1 U9849 ( .A(n3841), .B(n5415), .Z(N327) );
  CEOX1 U9850 ( .A(N326), .B(mem_data1[308]), .Z(N7971) );
  CNR2X1 U9851 ( .A(n3840), .B(n5414), .Z(N326) );
  CEOX1 U9852 ( .A(N325), .B(mem_data1[307]), .Z(N7972) );
  CNR2X1 U9853 ( .A(n3839), .B(n5413), .Z(N325) );
  CEOX1 U9854 ( .A(N324), .B(mem_data1[306]), .Z(N7973) );
  CNR2X1 U9855 ( .A(n3838), .B(n5412), .Z(N324) );
  CEOX1 U9856 ( .A(N320), .B(mem_data1[302]), .Z(N7977) );
  CNR2X1 U9857 ( .A(n3834), .B(n5408), .Z(N320) );
  CEOX1 U9858 ( .A(mem_data1[295]), .B(N313), .Z(N7984) );
  CNR2IX1 U9859 ( .B(n3831), .A(n5400), .Z(N313) );
  CEOX1 U9860 ( .A(N307), .B(mem_data1[289]), .Z(N7990) );
  CNR2X1 U9861 ( .A(n3845), .B(n5393), .Z(N307) );
  CEOX1 U9862 ( .A(N303), .B(mem_data1[285]), .Z(N7994) );
  CNR2X1 U9863 ( .A(n3841), .B(n5389), .Z(N303) );
  CEOX1 U9864 ( .A(N293), .B(mem_data1[275]), .Z(N8004) );
  CNR2X1 U9865 ( .A(n3838), .B(n5378), .Z(N293) );
  CEOX1 U9866 ( .A(N285), .B(mem_data1[267]), .Z(N8012) );
  CNR2X1 U9867 ( .A(n3847), .B(n5368), .Z(N285) );
  CEOX1 U9868 ( .A(N281), .B(mem_data1[263]), .Z(N8016) );
  CNR2X1 U9869 ( .A(n3844), .B(n5364), .Z(N281) );
  CEOX1 U9870 ( .A(N279), .B(mem_data1[261]), .Z(N8018) );
  CNR2X1 U9871 ( .A(n3842), .B(n5361), .Z(N279) );
  CEOX1 U9872 ( .A(N249), .B(mem_data1[231]), .Z(N8048) );
  CEOX1 U9873 ( .A(N247), .B(mem_data1[229]), .Z(N8050) );
  CEOX1 U9874 ( .A(N207), .B(mem_data1[189]), .Z(N8090) );
  CNR2X1 U9875 ( .A(n3830), .B(n5877), .Z(N207) );
  CEOX1 U9876 ( .A(N145), .B(mem_data1[127]), .Z(N8152) );
  CEOX1 U9877 ( .A(N115), .B(mem_data1[97]), .Z(N8182) );
  CEOX1 U9878 ( .A(N81), .B(mem_data1[63]), .Z(N8216) );
  CNR2X1 U9879 ( .A(n3841), .B(n5919), .Z(N81) );
  CEOX1 U9880 ( .A(N79), .B(mem_data1[61]), .Z(N8218) );
  CNR2X1 U9881 ( .A(n3845), .B(n5877), .Z(N79) );
  CEOX1 U9882 ( .A(N78), .B(mem_data1[60]), .Z(N8219) );
  CEOX1 U9883 ( .A(N1031), .B(mem_data1[1013]), .Z(N7266) );
  CNR2X1 U9884 ( .A(n3833), .B(n6371), .Z(N1031) );
  CEOX1 U9885 ( .A(N1030), .B(mem_data1[1012]), .Z(N7267) );
  CNR2X1 U9886 ( .A(n3817), .B(n6369), .Z(N1030) );
  CEOX1 U9887 ( .A(N1029), .B(mem_data1[1011]), .Z(N7268) );
  CNR2X1 U9888 ( .A(n3823), .B(n6367), .Z(N1029) );
  CEOX1 U9889 ( .A(N1028), .B(mem_data1[1010]), .Z(N7269) );
  CNR2X1 U9890 ( .A(n3821), .B(n6365), .Z(N1028) );
  CEOX1 U9891 ( .A(N1027), .B(mem_data1[1009]), .Z(N7270) );
  CNR2X1 U9892 ( .A(n3829), .B(n6363), .Z(N1027) );
  CEOX1 U9893 ( .A(N1026), .B(mem_data1[1008]), .Z(N7271) );
  CNR2X1 U9894 ( .A(n3820), .B(n6361), .Z(N1026) );
  CEOX1 U9895 ( .A(N1016), .B(mem_data1[998]), .Z(N7281) );
  CNR2X1 U9896 ( .A(n3824), .B(n6510), .Z(N1016) );
  CEOX1 U9897 ( .A(N670), .B(mem_data1[652]), .Z(N7627) );
  CNR2X1 U9898 ( .A(n3826), .B(n5933), .Z(N670) );
  CEOX1 U9899 ( .A(N542), .B(mem_data1[524]), .Z(N7755) );
  CNR2X1 U9900 ( .A(n3835), .B(n5933), .Z(N542) );
  CNR2IX1 U9901 ( .B(datain0[23]), .A(n4387), .Z(n5033) );
  CNR2IX1 U9902 ( .B(datain0[19]), .A(n4387), .Z(n5005) );
  CNR2IX1 U9903 ( .B(datain0[22]), .A(n4387), .Z(n5026) );
  CNR2IX1 U9904 ( .B(datain0[18]), .A(n4387), .Z(n4998) );
  CNR2IX1 U9905 ( .B(datain0[21]), .A(n4387), .Z(n5019) );
  CNR2IX1 U9906 ( .B(datain0[20]), .A(n4387), .Z(n5012) );
  CNR2IX1 U9907 ( .B(datain0[11]), .A(n4388), .Z(n4953) );
  CNR2IX1 U9908 ( .B(datain0[10]), .A(n4388), .Z(n4947) );
  CNR2IX1 U9909 ( .B(datain0[16]), .A(n4388), .Z(n4984) );
  CNR2IX1 U9910 ( .B(datain0[15]), .A(n4388), .Z(n4978) );
  CNR2IX1 U9911 ( .B(datain0[14]), .A(n4388), .Z(n4971) );
  CNR2IX1 U9912 ( .B(datain0[13]), .A(n4388), .Z(n4965) );
  CNR2IX1 U9913 ( .B(datain0[24]), .A(n4387), .Z(n5040) );
  CNR2IX1 U9914 ( .B(datain0[12]), .A(n4388), .Z(n4959) );
  CNR2IX1 U9915 ( .B(datain0[9]), .A(n4388), .Z(n4941) );
  CNR2IX1 U9916 ( .B(datain0[17]), .A(n4387), .Z(n4991) );
  COND1XL U9917 ( .A(n55), .B(n3238), .C(n56), .Z(n3173) );
  COND1XL U9918 ( .A(n55), .B(n3237), .C(n59), .Z(n3174) );
  COND1XL U9919 ( .A(n55), .B(n3236), .C(n60), .Z(n3175) );
  COND1XL U9920 ( .A(n55), .B(n3235), .C(n61), .Z(n3176) );
  COND1XL U9921 ( .A(n55), .B(n3234), .C(n62), .Z(n3177) );
  COND1XL U9922 ( .A(n55), .B(n3233), .C(n63), .Z(n3178) );
  COND1XL U9923 ( .A(n55), .B(n3232), .C(n64), .Z(n3179) );
  COND1XL U9924 ( .A(n55), .B(n3231), .C(n65), .Z(n3180) );
  COND1XL U9925 ( .A(n55), .B(n3230), .C(n66), .Z(n3181) );
  COND1XL U9926 ( .A(n55), .B(n3229), .C(n67), .Z(n3182) );
  COND1XL U9927 ( .A(n55), .B(n3228), .C(n68), .Z(n3183) );
  COND1XL U9928 ( .A(n55), .B(n3227), .C(n69), .Z(n3184) );
  COND1XL U9929 ( .A(n55), .B(n3226), .C(n70), .Z(n3185) );
  COND1XL U9930 ( .A(n55), .B(n3225), .C(n71), .Z(n3186) );
  COND1XL U9931 ( .A(n55), .B(n3224), .C(n72), .Z(n3187) );
  CND3XL U9932 ( .A(n632), .B(n633), .C(n634), .Z(N9814) );
  CND2X1 U9933 ( .A(N5648), .B(n3686), .Z(n633) );
  CND3XL U9934 ( .A(n635), .B(n636), .C(n637), .Z(N9813) );
  CND2X1 U9935 ( .A(N5647), .B(n3686), .Z(n636) );
  CND3XL U9936 ( .A(n638), .B(n639), .C(n640), .Z(N9812) );
  CND2X1 U9937 ( .A(N5646), .B(n3686), .Z(n639) );
  CND3XL U9938 ( .A(n644), .B(n645), .C(n646), .Z(N9810) );
  CND2X1 U9939 ( .A(N5644), .B(n3693), .Z(n645) );
  CND3XL U9940 ( .A(n647), .B(n648), .C(n649), .Z(N9809) );
  CND2X1 U9941 ( .A(N5643), .B(n3697), .Z(n648) );
  CND3XL U9942 ( .A(n650), .B(n651), .C(n652), .Z(N9808) );
  CND2X1 U9943 ( .A(N5642), .B(n3688), .Z(n651) );
  CND3XL U9944 ( .A(n653), .B(n654), .C(n655), .Z(N9807) );
  CND2X1 U9945 ( .A(N5641), .B(n3691), .Z(n654) );
  CND3XL U9946 ( .A(n659), .B(n660), .C(n661), .Z(N9805) );
  CND2X1 U9947 ( .A(N5639), .B(n3696), .Z(n660) );
  CND3XL U9948 ( .A(n662), .B(n663), .C(n664), .Z(N9804) );
  CANR2X1 U9949 ( .A(N2556), .B(n3570), .C(n3607), .D(N7799), .Z(n664) );
  CND2X1 U9950 ( .A(N5638), .B(n3685), .Z(n663) );
  CND3XL U9951 ( .A(n671), .B(n672), .C(n673), .Z(N9801) );
  CND2X1 U9952 ( .A(N5635), .B(n3685), .Z(n672) );
  CND3XL U9953 ( .A(n677), .B(n678), .C(n679), .Z(N9799) );
  CND3XL U9954 ( .A(n707), .B(n708), .C(n709), .Z(N9789) );
  CND2X1 U9955 ( .A(N5623), .B(n3687), .Z(n708) );
  CND3XL U9956 ( .A(n710), .B(n711), .C(n712), .Z(N9788) );
  CND3XL U9957 ( .A(n713), .B(n714), .C(n715), .Z(N9787) );
  CND2X1 U9958 ( .A(N5621), .B(n3688), .Z(n714) );
  CND3XL U9959 ( .A(n719), .B(n720), .C(n721), .Z(N9785) );
  CND3XL U9960 ( .A(n722), .B(n723), .C(n724), .Z(N9784) );
  CND3XL U9961 ( .A(n731), .B(n732), .C(n733), .Z(N9781) );
  CND3XL U9962 ( .A(n737), .B(n738), .C(n739), .Z(N9779) );
  CND2X1 U9963 ( .A(N5613), .B(n3688), .Z(n738) );
  CND3XL U9964 ( .A(n743), .B(n744), .C(n745), .Z(N9777) );
  CND2X1 U9965 ( .A(N5611), .B(n3698), .Z(n744) );
  CND3XL U9966 ( .A(n749), .B(n750), .C(n751), .Z(N9775) );
  CND3XL U9967 ( .A(n752), .B(n753), .C(n754), .Z(N9774) );
  CND3XL U9968 ( .A(n761), .B(n762), .C(n763), .Z(N9771) );
  CND3XL U9969 ( .A(n770), .B(n771), .C(n772), .Z(N9768) );
  CND2X1 U9970 ( .A(N5602), .B(n3686), .Z(n771) );
  CND3XL U9971 ( .A(n773), .B(n774), .C(n775), .Z(N9767) );
  CND3XL U9972 ( .A(n776), .B(n777), .C(n778), .Z(N9766) );
  CND2X1 U9973 ( .A(N5600), .B(n3688), .Z(n777) );
  CND3XL U9974 ( .A(n779), .B(n780), .C(n781), .Z(N9765) );
  CND2X1 U9975 ( .A(N5599), .B(n3690), .Z(n780) );
  CND3XL U9976 ( .A(n782), .B(n783), .C(n784), .Z(N9764) );
  CND2X1 U9977 ( .A(N5598), .B(n3683), .Z(n783) );
  CND3XL U9978 ( .A(n788), .B(n789), .C(n790), .Z(N9762) );
  CND2X1 U9979 ( .A(N5596), .B(n3689), .Z(n789) );
  CND3XL U9980 ( .A(n791), .B(n792), .C(n793), .Z(N9761) );
  CND2X1 U9981 ( .A(N5595), .B(n3693), .Z(n792) );
  CND3XL U9982 ( .A(n794), .B(n795), .C(n796), .Z(N9760) );
  CND2X1 U9983 ( .A(N5594), .B(n3688), .Z(n795) );
  CND3XL U9984 ( .A(n797), .B(n798), .C(n799), .Z(N9759) );
  CND2X1 U9985 ( .A(N5593), .B(n3697), .Z(n798) );
  CND3XL U9986 ( .A(n800), .B(n801), .C(n802), .Z(N9758) );
  CND3XL U9987 ( .A(n803), .B(n804), .C(n805), .Z(N9757) );
  CND2X1 U9988 ( .A(N5591), .B(n3692), .Z(n804) );
  CND3XL U9989 ( .A(n809), .B(n810), .C(n811), .Z(N9755) );
  CND2X1 U9990 ( .A(N5589), .B(n3685), .Z(n810) );
  CND3XL U9991 ( .A(n812), .B(n813), .C(n814), .Z(N9754) );
  CND2X1 U9992 ( .A(N5588), .B(n3684), .Z(n813) );
  CND3XL U9993 ( .A(n815), .B(n816), .C(n817), .Z(N9753) );
  CND3XL U9994 ( .A(n818), .B(n819), .C(n820), .Z(N9752) );
  CND2X1 U9995 ( .A(N5586), .B(n3691), .Z(n819) );
  CND3XL U9996 ( .A(n821), .B(n822), .C(n823), .Z(N9751) );
  CND2X1 U9997 ( .A(N5585), .B(n3684), .Z(n822) );
  CND3XL U9998 ( .A(n824), .B(n825), .C(n826), .Z(N9750) );
  CND2X1 U9999 ( .A(N5584), .B(n3693), .Z(n825) );
  CND3XL U10000 ( .A(n827), .B(n828), .C(n829), .Z(N9749) );
  CND2X1 U10001 ( .A(N5583), .B(n3695), .Z(n828) );
  CND3XL U10002 ( .A(n833), .B(n834), .C(n835), .Z(N9747) );
  CND2X1 U10003 ( .A(N5581), .B(n3691), .Z(n834) );
  CND3XL U10004 ( .A(n839), .B(n840), .C(n841), .Z(N9745) );
  CND2X1 U10005 ( .A(N5579), .B(n3695), .Z(n840) );
  CND3XL U10006 ( .A(n845), .B(n846), .C(n847), .Z(N9743) );
  CND2X1 U10007 ( .A(N5577), .B(n3689), .Z(n846) );
  CND3XL U10008 ( .A(n848), .B(n849), .C(n850), .Z(N9742) );
  CND3XL U10009 ( .A(n866), .B(n867), .C(n868), .Z(N9736) );
  CND3XL U10010 ( .A(n869), .B(n870), .C(n871), .Z(N9735) );
  CND3XL U10011 ( .A(n872), .B(n873), .C(n874), .Z(N9734) );
  CND3XL U10012 ( .A(n899), .B(n900), .C(n901), .Z(N9725) );
  CND2X1 U10013 ( .A(N5559), .B(n3689), .Z(n900) );
  CND3XL U10014 ( .A(n905), .B(n906), .C(n907), .Z(N9723) );
  CND2X1 U10015 ( .A(N5557), .B(n3686), .Z(n906) );
  CND3XL U10016 ( .A(n908), .B(n909), .C(n910), .Z(N9722) );
  CND3XL U10017 ( .A(n911), .B(n912), .C(n913), .Z(N9721) );
  CND3XL U10018 ( .A(n914), .B(n915), .C(n916), .Z(N9720) );
  CND3XL U10019 ( .A(n917), .B(n918), .C(n919), .Z(N9719) );
  CND2X1 U10020 ( .A(N5553), .B(n3690), .Z(n918) );
  CND3XL U10021 ( .A(n923), .B(n924), .C(n925), .Z(N9717) );
  CND3XL U10022 ( .A(n929), .B(n930), .C(n931), .Z(N9715) );
  CND2X1 U10023 ( .A(N5549), .B(n3685), .Z(n930) );
  CND3XL U10024 ( .A(n935), .B(n936), .C(n937), .Z(N9713) );
  CND3XL U10025 ( .A(n938), .B(n939), .C(n940), .Z(N9712) );
  CND3XL U10026 ( .A(n941), .B(n942), .C(n943), .Z(N9711) );
  CND3XL U10027 ( .A(n944), .B(n945), .C(n946), .Z(N9710) );
  CND3XL U10028 ( .A(n968), .B(n969), .C(n970), .Z(N9702) );
  CND2X1 U10029 ( .A(N5536), .B(n3684), .Z(n969) );
  CND3XL U10030 ( .A(n980), .B(n981), .C(n982), .Z(N9698) );
  CND2X1 U10031 ( .A(N5532), .B(n3687), .Z(n981) );
  CND3XL U10032 ( .A(n992), .B(n993), .C(n994), .Z(N9694) );
  CANR2X1 U10033 ( .A(N2446), .B(n3581), .C(n3616), .D(N7909), .Z(n994) );
  CND2X1 U10034 ( .A(N5528), .B(n3693), .Z(n993) );
  CND3XL U10035 ( .A(n995), .B(n996), .C(n997), .Z(N9693) );
  CND2X1 U10036 ( .A(N5527), .B(n3686), .Z(n996) );
  CND3XL U10037 ( .A(n1001), .B(n1002), .C(n1003), .Z(N9691) );
  CND2X1 U10038 ( .A(N5525), .B(n3690), .Z(n1002) );
  CND3XL U10039 ( .A(n1007), .B(n1008), .C(n1009), .Z(N9689) );
  CND2X1 U10040 ( .A(N5523), .B(n3687), .Z(n1008) );
  CND3XL U10041 ( .A(n1013), .B(n1014), .C(n1015), .Z(N9687) );
  CND2X1 U10042 ( .A(N5521), .B(n3696), .Z(n1014) );
  CND3XL U10043 ( .A(n1016), .B(n1017), .C(n1018), .Z(N9686) );
  CND2X1 U10044 ( .A(N5520), .B(n3694), .Z(n1017) );
  CND3XL U10045 ( .A(n1019), .B(n1020), .C(n1021), .Z(N9685) );
  CND2X1 U10046 ( .A(N5519), .B(n3695), .Z(n1020) );
  CND3XL U10047 ( .A(n1025), .B(n1026), .C(n1027), .Z(N9683) );
  CND2X1 U10048 ( .A(N5517), .B(n3689), .Z(n1026) );
  CND3XL U10049 ( .A(n1040), .B(n1041), .C(n1042), .Z(N9678) );
  CND2X1 U10050 ( .A(N5512), .B(n3691), .Z(n1041) );
  CND3XL U10051 ( .A(n1043), .B(n1044), .C(n1045), .Z(N9677) );
  CND2X1 U10052 ( .A(N5511), .B(n3690), .Z(n1044) );
  CND3XL U10053 ( .A(n1052), .B(n1053), .C(n1054), .Z(N9674) );
  CND3XL U10054 ( .A(n1055), .B(n1056), .C(n1057), .Z(N9673) );
  CND2X1 U10055 ( .A(N5507), .B(n3690), .Z(n1056) );
  CND3XL U10056 ( .A(n1058), .B(n1059), .C(n1060), .Z(N9672) );
  CND3XL U10057 ( .A(n1064), .B(n1065), .C(n1066), .Z(N9670) );
  CND3XL U10058 ( .A(n1067), .B(n1068), .C(n1069), .Z(N9669) );
  CND3XL U10059 ( .A(n1070), .B(n1071), .C(n1072), .Z(N9668) );
  CND3XL U10060 ( .A(n1073), .B(n1074), .C(n1075), .Z(N9667) );
  CND3XL U10061 ( .A(n1076), .B(n1077), .C(n1078), .Z(N9666) );
  CND3XL U10062 ( .A(n1079), .B(n1080), .C(n1081), .Z(N9665) );
  CND3XL U10063 ( .A(n1082), .B(n1083), .C(n1084), .Z(N9664) );
  CND3XL U10064 ( .A(n1085), .B(n1086), .C(n1087), .Z(N9663) );
  CND2X1 U10065 ( .A(N5497), .B(n3690), .Z(n1086) );
  CND3XL U10066 ( .A(n1091), .B(n1092), .C(n1093), .Z(N9661) );
  CND3XL U10067 ( .A(n1097), .B(n1098), .C(n1099), .Z(N9659) );
  CND2X1 U10068 ( .A(N5493), .B(n3696), .Z(n1098) );
  CND3XL U10069 ( .A(n1121), .B(n1122), .C(n1123), .Z(N9651) );
  CND2X1 U10070 ( .A(N5485), .B(n3687), .Z(n1122) );
  CND3XL U10071 ( .A(n1124), .B(n1125), .C(n1126), .Z(N9650) );
  CND3XL U10072 ( .A(n1127), .B(n1128), .C(n1129), .Z(N9649) );
  CND2X1 U10073 ( .A(N5483), .B(n3683), .Z(n1128) );
  CND3XL U10074 ( .A(n1130), .B(n1131), .C(n1132), .Z(N9648) );
  CND3XL U10075 ( .A(n1133), .B(n1134), .C(n1135), .Z(N9647) );
  CND3XL U10076 ( .A(n1139), .B(n1140), .C(n1141), .Z(N9645) );
  CND3XL U10077 ( .A(n1142), .B(n1143), .C(n1144), .Z(N9644) );
  CANR2X1 U10078 ( .A(N2396), .B(n3582), .C(n3617), .D(N7959), .Z(n1144) );
  CND2X1 U10079 ( .A(N5478), .B(n3683), .Z(n1143) );
  CND3XL U10080 ( .A(n1163), .B(n1164), .C(n1165), .Z(N9637) );
  CND2X1 U10081 ( .A(N5471), .B(n3684), .Z(n1164) );
  CND3XL U10082 ( .A(n1175), .B(n1176), .C(n1177), .Z(N9633) );
  CND2X1 U10083 ( .A(N5467), .B(n3691), .Z(n1176) );
  CND3XL U10084 ( .A(n1190), .B(n1191), .C(n1192), .Z(N9628) );
  CND3XL U10085 ( .A(n1199), .B(n1200), .C(n1201), .Z(N9625) );
  CND3XL U10086 ( .A(n1202), .B(n1203), .C(n1204), .Z(N9624) );
  CND2X1 U10087 ( .A(N5458), .B(n3690), .Z(n1203) );
  CND3XL U10088 ( .A(n1208), .B(n1209), .C(n1210), .Z(N9622) );
  CND2X1 U10089 ( .A(N5456), .B(n3698), .Z(n1209) );
  CND3XL U10090 ( .A(n1211), .B(n1212), .C(n1213), .Z(N9621) );
  CND2X1 U10091 ( .A(N5455), .B(n3698), .Z(n1212) );
  CND3XL U10092 ( .A(n1214), .B(n1215), .C(n1216), .Z(N9620) );
  CND2X1 U10093 ( .A(N5454), .B(n3689), .Z(n1215) );
  CND3XL U10094 ( .A(n1217), .B(n1218), .C(n1219), .Z(N9619) );
  CND2X1 U10095 ( .A(N5453), .B(n3689), .Z(n1218) );
  CND3XL U10096 ( .A(n1229), .B(n1230), .C(n1231), .Z(N9615) );
  CND2X1 U10097 ( .A(N5449), .B(n3686), .Z(n1230) );
  CND3XL U10098 ( .A(n1244), .B(n1245), .C(n1246), .Z(N9610) );
  CND3XL U10099 ( .A(n1253), .B(n1254), .C(n1255), .Z(N9607) );
  CND3XL U10100 ( .A(n1265), .B(n1266), .C(n1267), .Z(N9603) );
  CND3XL U10101 ( .A(n1268), .B(n1269), .C(n1270), .Z(N9602) );
  CND3XL U10102 ( .A(n1271), .B(n1272), .C(n1273), .Z(N9601) );
  CND3XL U10103 ( .A(n1283), .B(n1284), .C(n1285), .Z(N9597) );
  CND3XL U10104 ( .A(n1289), .B(n1290), .C(n1291), .Z(N9595) );
  CND2X1 U10105 ( .A(N5429), .B(n3683), .Z(n1290) );
  CND3XL U10106 ( .A(n1319), .B(n1320), .C(n1321), .Z(N9585) );
  CND2X1 U10107 ( .A(N5419), .B(n3689), .Z(n1320) );
  CND3XL U10108 ( .A(n1325), .B(n1326), .C(n1327), .Z(N9583) );
  CND3XL U10109 ( .A(n1331), .B(n1332), .C(n1333), .Z(N9581) );
  CND3XL U10110 ( .A(n1334), .B(n1335), .C(n1336), .Z(N9580) );
  CANR2X1 U10111 ( .A(N2332), .B(n3586), .C(n3621), .D(N8023), .Z(n1336) );
  CND2X1 U10112 ( .A(N5414), .B(n3694), .Z(n1335) );
  CND3XL U10113 ( .A(n1343), .B(n1344), .C(n1345), .Z(N9577) );
  CND2X1 U10114 ( .A(N5411), .B(n3695), .Z(n1344) );
  CND3XL U10115 ( .A(n1346), .B(n1347), .C(n1348), .Z(N9576) );
  CND2X1 U10116 ( .A(N5410), .B(n3688), .Z(n1347) );
  CND3XL U10117 ( .A(n1349), .B(n1350), .C(n1351), .Z(N9575) );
  CND2X1 U10118 ( .A(N5409), .B(n3693), .Z(n1350) );
  CND3XL U10119 ( .A(n1352), .B(n1353), .C(n1354), .Z(N9574) );
  CND2X1 U10120 ( .A(N5408), .B(n3691), .Z(n1353) );
  CND3XL U10121 ( .A(n1355), .B(n1356), .C(n1357), .Z(N9573) );
  CND2X1 U10122 ( .A(N5407), .B(n3686), .Z(n1356) );
  CND3XL U10123 ( .A(n1358), .B(n1359), .C(n1360), .Z(N9572) );
  CND2X1 U10124 ( .A(N5406), .B(n3693), .Z(n1359) );
  CND3XL U10125 ( .A(n1367), .B(n1368), .C(n1369), .Z(N9569) );
  CND2X1 U10126 ( .A(N5403), .B(n3683), .Z(n1368) );
  CND3XL U10127 ( .A(n1373), .B(n1374), .C(n1375), .Z(N9567) );
  CND2X1 U10128 ( .A(N5401), .B(n3690), .Z(n1374) );
  CND3XL U10129 ( .A(n1376), .B(n1377), .C(n1378), .Z(N9566) );
  CND3XL U10130 ( .A(n1442), .B(n1443), .C(n1444), .Z(N9544) );
  CND3XL U10131 ( .A(n1535), .B(n1536), .C(n1537), .Z(N9513) );
  CND2X1 U10132 ( .A(N5347), .B(n3694), .Z(n1536) );
  CND3XL U10133 ( .A(n1541), .B(n1542), .C(n1543), .Z(N9511) );
  CND3XL U10134 ( .A(n1544), .B(n1545), .C(n1546), .Z(N9510) );
  CND3XL U10135 ( .A(n1547), .B(n1548), .C(n1549), .Z(N9509) );
  CND3XL U10136 ( .A(n1553), .B(n1554), .C(n1555), .Z(N9507) );
  CND3XL U10137 ( .A(n1556), .B(n1557), .C(n1558), .Z(N9506) );
  CND3XL U10138 ( .A(n1559), .B(n1560), .C(n1561), .Z(N9505) );
  CND3XL U10139 ( .A(n1742), .B(n1743), .C(n1744), .Z(N9444) );
  CANR2X1 U10140 ( .A(N2196), .B(n3589), .C(n3623), .D(N8159), .Z(n1744) );
  CND2X1 U10141 ( .A(N5278), .B(n3697), .Z(n1743) );
  CND3XL U10142 ( .A(n1748), .B(n1749), .C(n1750), .Z(N9442) );
  CND2X1 U10143 ( .A(N5276), .B(n3697), .Z(n1749) );
  CND3XL U10144 ( .A(n1754), .B(n1755), .C(n1756), .Z(N9440) );
  CND2X1 U10145 ( .A(N5274), .B(n3697), .Z(n1755) );
  CND3XL U10146 ( .A(n1763), .B(n1764), .C(n1765), .Z(N9437) );
  CND3XL U10147 ( .A(n1769), .B(n1770), .C(n1771), .Z(N9435) );
  CND3XL U10148 ( .A(n1919), .B(n1920), .C(n1921), .Z(N9385) );
  CND2X1 U10149 ( .A(N5219), .B(n3684), .Z(n1920) );
  CND3XL U10150 ( .A(n1925), .B(n1926), .C(n1927), .Z(N9383) );
  CND3XL U10151 ( .A(n1928), .B(n1929), .C(n1930), .Z(N9382) );
  CNR2IX1 U10152 ( .B(datain0[7]), .A(n4389), .Z(n6056) );
  CAN2X1 U10153 ( .A(datain0[24]), .B(n4388), .Z(n5604) );
  CND3XL U10154 ( .A(n974), .B(n975), .C(n976), .Z(N9700) );
  CND2X1 U10155 ( .A(N5534), .B(n3689), .Z(n975) );
  CND3XL U10156 ( .A(n1061), .B(n1062), .C(n1063), .Z(N9671) );
  CND3XL U10157 ( .A(n2180), .B(n2181), .C(n2182), .Z(N10329) );
  CND3XL U10158 ( .A(n2183), .B(n2184), .C(n2185), .Z(N10328) );
  CND3XL U10159 ( .A(n2186), .B(n2187), .C(n2188), .Z(N10327) );
  CANR2X1 U10160 ( .A(N3079), .B(n3593), .C(n3627), .D(N7276), .Z(n2188) );
  CND2X1 U10161 ( .A(N6161), .B(n3689), .Z(n2187) );
  CANR2X1 U10162 ( .A(mem_data1[1003]), .B(n3898), .C(N9283), .D(n3673), .Z(
        n2186) );
  CND3XL U10163 ( .A(n2189), .B(n2190), .C(n2191), .Z(N10326) );
  CANR2X1 U10164 ( .A(N3078), .B(n3593), .C(n3627), .D(N7277), .Z(n2191) );
  CND2X1 U10165 ( .A(N6160), .B(n3693), .Z(n2190) );
  CANR2X1 U10166 ( .A(mem_data1[1002]), .B(n3898), .C(N9282), .D(n3673), .Z(
        n2189) );
  CND3XL U10167 ( .A(n2192), .B(n2193), .C(n2194), .Z(N10325) );
  CANR2X1 U10168 ( .A(N3077), .B(n3595), .C(n3627), .D(N7278), .Z(n2194) );
  CND2X1 U10169 ( .A(N6159), .B(n3690), .Z(n2193) );
  CANR2X1 U10170 ( .A(mem_data1[1001]), .B(n3898), .C(N9281), .D(n3673), .Z(
        n2192) );
  CND3XL U10171 ( .A(n2195), .B(n2196), .C(n2197), .Z(N10324) );
  CANR2X1 U10172 ( .A(N3076), .B(n3595), .C(n3627), .D(N7279), .Z(n2197) );
  CND2X1 U10173 ( .A(N6158), .B(n3685), .Z(n2196) );
  CANR2X1 U10174 ( .A(mem_data1[1000]), .B(n3898), .C(N9280), .D(n3673), .Z(
        n2195) );
  CND3XL U10175 ( .A(n2198), .B(n2199), .C(n2200), .Z(N10323) );
  CANR2X1 U10176 ( .A(N3075), .B(n3595), .C(n3629), .D(N7280), .Z(n2200) );
  CND2X1 U10177 ( .A(N6157), .B(n3694), .Z(n2199) );
  CANR2X1 U10178 ( .A(mem_data1[999]), .B(n3898), .C(N9279), .D(n3673), .Z(
        n2198) );
  CND3XL U10179 ( .A(n2201), .B(n2202), .C(n2203), .Z(N10322) );
  CANR2X1 U10180 ( .A(N3074), .B(n3595), .C(n3629), .D(N7281), .Z(n2203) );
  CND2X1 U10181 ( .A(N6156), .B(n3691), .Z(n2202) );
  CANR2X1 U10182 ( .A(mem_data1[998]), .B(n3898), .C(N9278), .D(n3673), .Z(
        n2201) );
  CND3XL U10183 ( .A(n2204), .B(n2205), .C(n2206), .Z(N10321) );
  CANR2X1 U10184 ( .A(N3073), .B(n3595), .C(n3629), .D(N7282), .Z(n2206) );
  CND2X1 U10185 ( .A(N6155), .B(n3694), .Z(n2205) );
  CANR2X1 U10186 ( .A(mem_data1[997]), .B(n3898), .C(N9277), .D(n3673), .Z(
        n2204) );
  CND3XL U10187 ( .A(n2207), .B(n2208), .C(n2209), .Z(N10320) );
  CANR2X1 U10188 ( .A(N3072), .B(n3595), .C(n3629), .D(N7283), .Z(n2209) );
  CND2X1 U10189 ( .A(N6154), .B(n3693), .Z(n2208) );
  CANR2X1 U10190 ( .A(mem_data1[996]), .B(n3898), .C(N9276), .D(n3673), .Z(
        n2207) );
  CND3XL U10191 ( .A(n2210), .B(n2211), .C(n2212), .Z(N10319) );
  CANR2X1 U10192 ( .A(N3071), .B(n3595), .C(n3629), .D(N7284), .Z(n2212) );
  CND2X1 U10193 ( .A(N6153), .B(n3693), .Z(n2211) );
  CANR2X1 U10194 ( .A(mem_data1[995]), .B(n3898), .C(N9275), .D(n3673), .Z(
        n2210) );
  CND3XL U10195 ( .A(n2213), .B(n2214), .C(n2215), .Z(N10318) );
  CANR2X1 U10196 ( .A(N3070), .B(n3595), .C(n3629), .D(N7285), .Z(n2215) );
  CND2X1 U10197 ( .A(N6152), .B(n3693), .Z(n2214) );
  CANR2X1 U10198 ( .A(mem_data1[994]), .B(n3898), .C(N9274), .D(n3673), .Z(
        n2213) );
  CND3XL U10199 ( .A(n2216), .B(n2217), .C(n2218), .Z(N10317) );
  CANR2X1 U10200 ( .A(N3069), .B(n3595), .C(n3629), .D(N7286), .Z(n2218) );
  CND2X1 U10201 ( .A(N6151), .B(n3693), .Z(n2217) );
  CANR2X1 U10202 ( .A(mem_data1[993]), .B(n3898), .C(N9273), .D(n3673), .Z(
        n2216) );
  CND3XL U10203 ( .A(n2219), .B(n2220), .C(n2221), .Z(N10316) );
  CANR2X1 U10204 ( .A(N3068), .B(n3595), .C(n3629), .D(N7287), .Z(n2221) );
  CND2X1 U10205 ( .A(N6150), .B(n3693), .Z(n2220) );
  CANR2X1 U10206 ( .A(mem_data1[992]), .B(n3898), .C(N9272), .D(n3673), .Z(
        n2219) );
  CND3XL U10207 ( .A(n2222), .B(n2223), .C(n2224), .Z(N10315) );
  CANR2X1 U10208 ( .A(N3067), .B(n3595), .C(n3629), .D(N7288), .Z(n2224) );
  CND2X1 U10209 ( .A(N6149), .B(n3693), .Z(n2223) );
  CANR2X1 U10210 ( .A(mem_data1[991]), .B(n3898), .C(N9271), .D(n3673), .Z(
        n2222) );
  CND3XL U10211 ( .A(n2225), .B(n2226), .C(n2227), .Z(N10314) );
  CANR2X1 U10212 ( .A(N3066), .B(n3595), .C(n3629), .D(N7289), .Z(n2227) );
  CND2X1 U10213 ( .A(N6148), .B(n3693), .Z(n2226) );
  CANR2X1 U10214 ( .A(mem_data1[990]), .B(n3898), .C(N9270), .D(n3673), .Z(
        n2225) );
  CND3XL U10215 ( .A(n2228), .B(n2229), .C(n2230), .Z(N10313) );
  CND3XL U10216 ( .A(n2231), .B(n2232), .C(n2233), .Z(N10312) );
  CND3XL U10217 ( .A(n2234), .B(n2235), .C(n2236), .Z(N10311) );
  CND3XL U10218 ( .A(n2237), .B(n2238), .C(n2239), .Z(N10310) );
  CND3XL U10219 ( .A(n2240), .B(n2241), .C(n2242), .Z(N10309) );
  CND3XL U10220 ( .A(n2243), .B(n2244), .C(n2245), .Z(N10308) );
  CND2X1 U10221 ( .A(N6142), .B(n3693), .Z(n2244) );
  CND3XL U10222 ( .A(n2246), .B(n2247), .C(n2248), .Z(N10307) );
  CND2X1 U10223 ( .A(N6141), .B(n3693), .Z(n2247) );
  CND3XL U10224 ( .A(n2249), .B(n2250), .C(n2251), .Z(N10306) );
  CND2X1 U10225 ( .A(N6140), .B(n3693), .Z(n2250) );
  CND3XL U10226 ( .A(n2252), .B(n2253), .C(n2254), .Z(N10305) );
  CANR2X1 U10227 ( .A(N3057), .B(n3594), .C(n3628), .D(N7298), .Z(n2254) );
  CND2X1 U10228 ( .A(N6139), .B(n3684), .Z(n2253) );
  CANR2X1 U10229 ( .A(mem_data1[981]), .B(n3898), .C(N9261), .D(n3672), .Z(
        n2252) );
  CND3XL U10230 ( .A(n2255), .B(n2256), .C(n2257), .Z(N10304) );
  CANR2X1 U10231 ( .A(N3056), .B(n3594), .C(n3628), .D(N7299), .Z(n2257) );
  CND2X1 U10232 ( .A(N6138), .B(n3684), .Z(n2256) );
  CANR2X1 U10233 ( .A(mem_data1[980]), .B(n3898), .C(N9260), .D(n3672), .Z(
        n2255) );
  CND3XL U10234 ( .A(n2258), .B(n2259), .C(n2260), .Z(N10303) );
  CANR2X1 U10235 ( .A(N3055), .B(n3594), .C(n3628), .D(N7300), .Z(n2260) );
  CND2X1 U10236 ( .A(N6137), .B(n3684), .Z(n2259) );
  CANR2X1 U10237 ( .A(mem_data1[979]), .B(n3898), .C(N9259), .D(n3672), .Z(
        n2258) );
  CND3XL U10238 ( .A(n2261), .B(n2262), .C(n2263), .Z(N10302) );
  CANR2X1 U10239 ( .A(N3054), .B(n3594), .C(n3628), .D(N7301), .Z(n2263) );
  CND2X1 U10240 ( .A(N6136), .B(n3684), .Z(n2262) );
  CANR2X1 U10241 ( .A(mem_data1[978]), .B(n3898), .C(N9258), .D(n3672), .Z(
        n2261) );
  CND3XL U10242 ( .A(n2264), .B(n2265), .C(n2266), .Z(N10301) );
  CANR2X1 U10243 ( .A(N3053), .B(n3596), .C(n3628), .D(N7302), .Z(n2266) );
  CND2X1 U10244 ( .A(N6135), .B(n3684), .Z(n2265) );
  CANR2X1 U10245 ( .A(mem_data1[977]), .B(n3898), .C(N9257), .D(n3672), .Z(
        n2264) );
  CND3XL U10246 ( .A(n2267), .B(n2268), .C(n2269), .Z(N10300) );
  CANR2X1 U10247 ( .A(N3052), .B(n3596), .C(n3628), .D(N7303), .Z(n2269) );
  CND2X1 U10248 ( .A(N6134), .B(n3684), .Z(n2268) );
  CANR2X1 U10249 ( .A(mem_data1[976]), .B(n3898), .C(N9256), .D(n3672), .Z(
        n2267) );
  CND3XL U10250 ( .A(n2270), .B(n2271), .C(n2272), .Z(N10299) );
  CANR2X1 U10251 ( .A(N3051), .B(n3596), .C(n3628), .D(N7304), .Z(n2272) );
  CND2X1 U10252 ( .A(N6133), .B(n3684), .Z(n2271) );
  CANR2X1 U10253 ( .A(mem_data1[975]), .B(n3898), .C(N9255), .D(n3672), .Z(
        n2270) );
  CND3XL U10254 ( .A(n2273), .B(n2274), .C(n2275), .Z(N10298) );
  CANR2X1 U10255 ( .A(N3050), .B(n3596), .C(n3628), .D(N7305), .Z(n2275) );
  CND2X1 U10256 ( .A(N6132), .B(n3684), .Z(n2274) );
  CANR2X1 U10257 ( .A(mem_data1[974]), .B(n3898), .C(N9254), .D(n3672), .Z(
        n2273) );
  CND3XL U10258 ( .A(n2276), .B(n2277), .C(n2278), .Z(N10297) );
  CANR2X1 U10259 ( .A(N3049), .B(n3596), .C(n3630), .D(N7306), .Z(n2278) );
  CND2X1 U10260 ( .A(N6131), .B(n3684), .Z(n2277) );
  CANR2X1 U10261 ( .A(mem_data1[973]), .B(n3898), .C(N9253), .D(n3672), .Z(
        n2276) );
  CND3XL U10262 ( .A(n2279), .B(n2280), .C(n2281), .Z(N10296) );
  CANR2X1 U10263 ( .A(N3048), .B(n3596), .C(n3630), .D(N7307), .Z(n2281) );
  CND2X1 U10264 ( .A(N6130), .B(n3684), .Z(n2280) );
  CANR2X1 U10265 ( .A(mem_data1[972]), .B(n3898), .C(N9252), .D(n3672), .Z(
        n2279) );
  CND3XL U10266 ( .A(n2282), .B(n2283), .C(n2284), .Z(N10295) );
  CANR2X1 U10267 ( .A(N3047), .B(n3596), .C(n3630), .D(N7308), .Z(n2284) );
  CND2X1 U10268 ( .A(N6129), .B(n3695), .Z(n2283) );
  CANR2X1 U10269 ( .A(mem_data1[971]), .B(n3898), .C(N9251), .D(n3672), .Z(
        n2282) );
  CND3XL U10270 ( .A(n2285), .B(n2286), .C(n2287), .Z(N10294) );
  CANR2X1 U10271 ( .A(N3046), .B(n3596), .C(n3630), .D(N7309), .Z(n2287) );
  CND2X1 U10272 ( .A(N6128), .B(n3690), .Z(n2286) );
  CANR2X1 U10273 ( .A(mem_data1[970]), .B(n3898), .C(N9250), .D(n3672), .Z(
        n2285) );
  CND3XL U10274 ( .A(n2288), .B(n2289), .C(n2290), .Z(N10293) );
  CANR2X1 U10275 ( .A(N3045), .B(n3596), .C(n3630), .D(N7310), .Z(n2290) );
  CND2X1 U10276 ( .A(N6127), .B(n3685), .Z(n2289) );
  CANR2X1 U10277 ( .A(mem_data1[969]), .B(n3898), .C(N9249), .D(n3672), .Z(
        n2288) );
  CND3XL U10278 ( .A(n2291), .B(n2292), .C(n2293), .Z(N10292) );
  CANR2X1 U10279 ( .A(N3044), .B(n3596), .C(n3630), .D(N7311), .Z(n2293) );
  CND2X1 U10280 ( .A(N6126), .B(n3695), .Z(n2292) );
  CANR2X1 U10281 ( .A(mem_data1[968]), .B(n3898), .C(N9248), .D(n3672), .Z(
        n2291) );
  CND3XL U10282 ( .A(n2294), .B(n2295), .C(n2296), .Z(N10291) );
  CANR2X1 U10283 ( .A(N3043), .B(n3596), .C(n3630), .D(N7312), .Z(n2296) );
  CND2X1 U10284 ( .A(N6125), .B(n3695), .Z(n2295) );
  CANR2X1 U10285 ( .A(mem_data1[967]), .B(n3898), .C(N9247), .D(n3672), .Z(
        n2294) );
  CND3XL U10286 ( .A(n2297), .B(n2298), .C(n2299), .Z(N10290) );
  CANR2X1 U10287 ( .A(N3042), .B(n3596), .C(n3630), .D(N7313), .Z(n2299) );
  CND2X1 U10288 ( .A(N6124), .B(n3696), .Z(n2298) );
  CANR2X1 U10289 ( .A(mem_data1[966]), .B(n3898), .C(N9246), .D(n3672), .Z(
        n2297) );
  CND3XL U10290 ( .A(n2300), .B(n2301), .C(n2302), .Z(N10289) );
  CANR2X1 U10291 ( .A(N3041), .B(n3596), .C(n3630), .D(N7314), .Z(n2302) );
  CND2X1 U10292 ( .A(N6123), .B(n3688), .Z(n2301) );
  CANR2X1 U10293 ( .A(mem_data1[965]), .B(n3898), .C(N9245), .D(n3672), .Z(
        n2300) );
  CND3XL U10294 ( .A(n2303), .B(n2304), .C(n2305), .Z(N10288) );
  CANR2X1 U10295 ( .A(N3040), .B(n3596), .C(n3630), .D(N7315), .Z(n2305) );
  CND2X1 U10296 ( .A(N6122), .B(n3686), .Z(n2304) );
  CANR2X1 U10297 ( .A(mem_data1[964]), .B(n3898), .C(N9244), .D(n3672), .Z(
        n2303) );
  CND3XL U10298 ( .A(n2306), .B(n2307), .C(n2308), .Z(N10287) );
  CANR2X1 U10299 ( .A(N3039), .B(n3595), .C(n3630), .D(N7316), .Z(n2308) );
  CND2X1 U10300 ( .A(N6121), .B(n3687), .Z(n2307) );
  CANR2X1 U10301 ( .A(mem_data1[963]), .B(n3898), .C(N9243), .D(n3672), .Z(
        n2306) );
  CND3XL U10302 ( .A(n2309), .B(n2310), .C(n2311), .Z(N10286) );
  CANR2X1 U10303 ( .A(N3038), .B(n3595), .C(n3630), .D(N7317), .Z(n2311) );
  CND2X1 U10304 ( .A(N6120), .B(n3696), .Z(n2310) );
  CANR2X1 U10305 ( .A(mem_data1[962]), .B(n3898), .C(N9242), .D(n3672), .Z(
        n2309) );
  CND3XL U10306 ( .A(n2312), .B(n2313), .C(n2314), .Z(N10285) );
  CANR2X1 U10307 ( .A(N3037), .B(n3595), .C(n3629), .D(N7318), .Z(n2314) );
  CND2X1 U10308 ( .A(N6119), .B(n3698), .Z(n2313) );
  CANR2X1 U10309 ( .A(mem_data1[961]), .B(n3898), .C(N9241), .D(n3673), .Z(
        n2312) );
  CND3XL U10310 ( .A(n2315), .B(n2316), .C(n2317), .Z(N10284) );
  CANR2X1 U10311 ( .A(N3036), .B(n3595), .C(n3629), .D(N7319), .Z(n2317) );
  CND2X1 U10312 ( .A(N6118), .B(n3684), .Z(n2316) );
  CANR2X1 U10313 ( .A(mem_data1[960]), .B(n3898), .C(N9240), .D(n3673), .Z(
        n2315) );
  CND3XL U10314 ( .A(n2318), .B(n2319), .C(n2320), .Z(N10283) );
  CANR2X1 U10315 ( .A(N3035), .B(n3595), .C(n3629), .D(N7320), .Z(n2320) );
  CND2X1 U10316 ( .A(N6117), .B(n3686), .Z(n2319) );
  CANR2X1 U10317 ( .A(mem_data1[959]), .B(n3898), .C(N9239), .D(n3671), .Z(
        n2318) );
  CND3XL U10318 ( .A(n2321), .B(n2322), .C(n2323), .Z(N10282) );
  CANR2X1 U10319 ( .A(N3034), .B(n3595), .C(n3629), .D(N7321), .Z(n2323) );
  CND2X1 U10320 ( .A(N6116), .B(n3693), .Z(n2322) );
  CANR2X1 U10321 ( .A(mem_data1[958]), .B(n3898), .C(N9238), .D(n3671), .Z(
        n2321) );
  CND3XL U10322 ( .A(n2324), .B(n2325), .C(n2326), .Z(N10281) );
  CND3XL U10323 ( .A(n2327), .B(n2328), .C(n2329), .Z(N10280) );
  CANR2X1 U10324 ( .A(N3032), .B(n3595), .C(n3629), .D(N7323), .Z(n2329) );
  CND2X1 U10325 ( .A(N6114), .B(n3683), .Z(n2328) );
  CANR2X1 U10326 ( .A(mem_data1[956]), .B(n3898), .C(N9236), .D(n3671), .Z(
        n2327) );
  CND3XL U10327 ( .A(n2330), .B(n2331), .C(n2332), .Z(N10279) );
  CANR2X1 U10328 ( .A(N3031), .B(n3595), .C(n3629), .D(N7324), .Z(n2332) );
  CND2X1 U10329 ( .A(N6113), .B(n3685), .Z(n2331) );
  CANR2X1 U10330 ( .A(mem_data1[955]), .B(n3898), .C(N9235), .D(n3671), .Z(
        n2330) );
  CND3XL U10331 ( .A(n2333), .B(n2334), .C(n2335), .Z(N10278) );
  CANR2X1 U10332 ( .A(N3030), .B(n3595), .C(n3629), .D(N7325), .Z(n2335) );
  CND2X1 U10333 ( .A(N6112), .B(n3697), .Z(n2334) );
  CANR2X1 U10334 ( .A(mem_data1[954]), .B(n3898), .C(N9234), .D(n3671), .Z(
        n2333) );
  CND3XL U10335 ( .A(n2336), .B(n2337), .C(n2338), .Z(N10277) );
  CANR2X1 U10336 ( .A(N3029), .B(n3595), .C(n3629), .D(N7326), .Z(n2338) );
  CND2X1 U10337 ( .A(N6111), .B(n3691), .Z(n2337) );
  CANR2X1 U10338 ( .A(mem_data1[953]), .B(n3898), .C(N9233), .D(n3671), .Z(
        n2336) );
  CND3XL U10339 ( .A(n2339), .B(n2340), .C(n2341), .Z(N10276) );
  CANR2X1 U10340 ( .A(N3028), .B(n3588), .C(n3629), .D(N7327), .Z(n2341) );
  CND2X1 U10341 ( .A(N6110), .B(n3694), .Z(n2340) );
  CANR2X1 U10342 ( .A(mem_data1[952]), .B(n3898), .C(N9232), .D(n3671), .Z(
        n2339) );
  CND3XL U10343 ( .A(n2342), .B(n2343), .C(n2344), .Z(N10275) );
  CANR2X1 U10344 ( .A(N3027), .B(n3588), .C(n3629), .D(N7328), .Z(n2344) );
  CND2X1 U10345 ( .A(N6109), .B(n3689), .Z(n2343) );
  CANR2X1 U10346 ( .A(mem_data1[951]), .B(n3898), .C(N9231), .D(n3671), .Z(
        n2342) );
  CND3XL U10347 ( .A(n2345), .B(n2346), .C(n2347), .Z(N10274) );
  CANR2X1 U10348 ( .A(N3026), .B(n3588), .C(n3629), .D(N7329), .Z(n2347) );
  CND2X1 U10349 ( .A(N6108), .B(n3688), .Z(n2346) );
  CANR2X1 U10350 ( .A(mem_data1[950]), .B(n3898), .C(N9230), .D(n3671), .Z(
        n2345) );
  CND3XL U10351 ( .A(n2348), .B(n2349), .C(n2350), .Z(N10273) );
  CANR2X1 U10352 ( .A(N3025), .B(n3588), .C(n3629), .D(N7330), .Z(n2350) );
  CND2X1 U10353 ( .A(N6107), .B(n3684), .Z(n2349) );
  CANR2X1 U10354 ( .A(mem_data1[949]), .B(n3898), .C(N9229), .D(n3671), .Z(
        n2348) );
  CND3XL U10355 ( .A(n2351), .B(n2352), .C(n2353), .Z(N10272) );
  CANR2X1 U10356 ( .A(N3024), .B(n3588), .C(n3629), .D(N7331), .Z(n2353) );
  CND2X1 U10357 ( .A(N6106), .B(n3684), .Z(n2352) );
  CANR2X1 U10358 ( .A(mem_data1[948]), .B(n3898), .C(N9228), .D(n3671), .Z(
        n2351) );
  CND3XL U10359 ( .A(n2354), .B(n2355), .C(n2356), .Z(N10271) );
  CANR2X1 U10360 ( .A(N3023), .B(n3588), .C(n3629), .D(N7332), .Z(n2356) );
  CND2X1 U10361 ( .A(N6105), .B(n3684), .Z(n2355) );
  CANR2X1 U10362 ( .A(mem_data1[947]), .B(n3898), .C(N9227), .D(n3671), .Z(
        n2354) );
  CND3XL U10363 ( .A(n2357), .B(n2358), .C(n2359), .Z(N10270) );
  CANR2X1 U10364 ( .A(N3022), .B(n3588), .C(n3622), .D(N7333), .Z(n2359) );
  CND2X1 U10365 ( .A(N6104), .B(n3684), .Z(n2358) );
  CANR2X1 U10366 ( .A(mem_data1[946]), .B(n3898), .C(N9226), .D(n3671), .Z(
        n2357) );
  CND3XL U10367 ( .A(n2360), .B(n2361), .C(n2362), .Z(N10269) );
  CANR2X1 U10368 ( .A(N3021), .B(n3587), .C(n3622), .D(N7334), .Z(n2362) );
  CND2X1 U10369 ( .A(N6103), .B(n3684), .Z(n2361) );
  CANR2X1 U10370 ( .A(mem_data1[945]), .B(n3898), .C(N9225), .D(n3671), .Z(
        n2360) );
  CND3XL U10371 ( .A(n2363), .B(n2364), .C(n2365), .Z(N10268) );
  CANR2X1 U10372 ( .A(N3020), .B(n3587), .C(n3622), .D(N7335), .Z(n2365) );
  CND2X1 U10373 ( .A(N6102), .B(n3684), .Z(n2364) );
  CANR2X1 U10374 ( .A(mem_data1[944]), .B(n3898), .C(N9224), .D(n3671), .Z(
        n2363) );
  CND3XL U10375 ( .A(n2366), .B(n2367), .C(n2368), .Z(N10267) );
  CANR2X1 U10376 ( .A(N3019), .B(n3587), .C(n3622), .D(N7336), .Z(n2368) );
  CND2X1 U10377 ( .A(N6101), .B(n3684), .Z(n2367) );
  CANR2X1 U10378 ( .A(mem_data1[943]), .B(n3898), .C(N9223), .D(n3671), .Z(
        n2366) );
  CND3XL U10379 ( .A(n2369), .B(n2370), .C(n2371), .Z(N10266) );
  CANR2X1 U10380 ( .A(N3018), .B(n3587), .C(n3622), .D(N7337), .Z(n2371) );
  CND2X1 U10381 ( .A(N6100), .B(n3684), .Z(n2370) );
  CANR2X1 U10382 ( .A(mem_data1[942]), .B(n3898), .C(N9222), .D(n3671), .Z(
        n2369) );
  CND3XL U10383 ( .A(n2372), .B(n2373), .C(n2374), .Z(N10265) );
  CANR2X1 U10384 ( .A(N3017), .B(n3587), .C(n3622), .D(N7338), .Z(n2374) );
  CND2X1 U10385 ( .A(N6099), .B(n3684), .Z(n2373) );
  CANR2X1 U10386 ( .A(mem_data1[941]), .B(n3898), .C(N9221), .D(n3671), .Z(
        n2372) );
  CND3XL U10387 ( .A(n2375), .B(n2376), .C(n2377), .Z(N10264) );
  CANR2X1 U10388 ( .A(N3016), .B(n3587), .C(n3622), .D(N7339), .Z(n2377) );
  CND2X1 U10389 ( .A(N6098), .B(n3684), .Z(n2376) );
  CANR2X1 U10390 ( .A(mem_data1[940]), .B(n3898), .C(N9220), .D(n3671), .Z(
        n2375) );
  CND3XL U10391 ( .A(n2378), .B(n2379), .C(n2380), .Z(N10263) );
  CANR2X1 U10392 ( .A(N3015), .B(n3587), .C(n3622), .D(N7340), .Z(n2380) );
  CND2X1 U10393 ( .A(N6097), .B(n3684), .Z(n2379) );
  CANR2X1 U10394 ( .A(mem_data1[939]), .B(n3898), .C(N9219), .D(n3671), .Z(
        n2378) );
  CND3XL U10395 ( .A(n2381), .B(n2382), .C(n2383), .Z(N10262) );
  CANR2X1 U10396 ( .A(N3014), .B(n3587), .C(n3622), .D(N7341), .Z(n2383) );
  CND2X1 U10397 ( .A(N6096), .B(n3684), .Z(n2382) );
  CANR2X1 U10398 ( .A(mem_data1[938]), .B(n3898), .C(N9218), .D(n3671), .Z(
        n2381) );
  CND3XL U10399 ( .A(n2384), .B(n2385), .C(n2386), .Z(N10261) );
  CANR2X1 U10400 ( .A(N3013), .B(n3589), .C(n3622), .D(N7342), .Z(n2386) );
  CND2X1 U10401 ( .A(N6095), .B(n3689), .Z(n2385) );
  CANR2X1 U10402 ( .A(mem_data1[937]), .B(n3898), .C(N9217), .D(n3670), .Z(
        n2384) );
  CND3XL U10403 ( .A(n2387), .B(n2388), .C(n2389), .Z(N10260) );
  CANR2X1 U10404 ( .A(N3012), .B(n3596), .C(n3622), .D(N7343), .Z(n2389) );
  CND2X1 U10405 ( .A(N6094), .B(n3695), .Z(n2388) );
  CANR2X1 U10406 ( .A(mem_data1[936]), .B(n3898), .C(N9216), .D(n3670), .Z(
        n2387) );
  CND3XL U10407 ( .A(n2390), .B(n2391), .C(n2392), .Z(N10259) );
  CANR2X1 U10408 ( .A(N3011), .B(n3595), .C(n3629), .D(N7344), .Z(n2392) );
  CND2X1 U10409 ( .A(N6093), .B(n3683), .Z(n2391) );
  CANR2X1 U10410 ( .A(mem_data1[935]), .B(n3898), .C(N9215), .D(n3670), .Z(
        n2390) );
  CND3XL U10411 ( .A(n2393), .B(n2394), .C(n2395), .Z(N10258) );
  CANR2X1 U10412 ( .A(N3010), .B(n3600), .C(n3632), .D(N7345), .Z(n2395) );
  CND2X1 U10413 ( .A(N6092), .B(n3693), .Z(n2394) );
  CANR2X1 U10414 ( .A(mem_data1[934]), .B(n3898), .C(N9214), .D(n3670), .Z(
        n2393) );
  CND3XL U10415 ( .A(n2396), .B(n2397), .C(n2398), .Z(N10257) );
  CANR2X1 U10416 ( .A(N3009), .B(n3600), .C(n3634), .D(N7346), .Z(n2398) );
  CND2X1 U10417 ( .A(N6091), .B(n3683), .Z(n2397) );
  CANR2X1 U10418 ( .A(mem_data1[933]), .B(n3898), .C(N9213), .D(n3670), .Z(
        n2396) );
  CND3XL U10419 ( .A(n2399), .B(n2400), .C(n2401), .Z(N10256) );
  CANR2X1 U10420 ( .A(N3008), .B(n3600), .C(n3634), .D(N7347), .Z(n2401) );
  CND2X1 U10421 ( .A(N6090), .B(n3688), .Z(n2400) );
  CANR2X1 U10422 ( .A(mem_data1[932]), .B(n3898), .C(N9212), .D(n3670), .Z(
        n2399) );
  CND3XL U10423 ( .A(n2402), .B(n2403), .C(n2404), .Z(N10255) );
  CANR2X1 U10424 ( .A(N3007), .B(n3600), .C(n3634), .D(N7348), .Z(n2404) );
  CND2X1 U10425 ( .A(N6089), .B(n3689), .Z(n2403) );
  CANR2X1 U10426 ( .A(mem_data1[931]), .B(n3898), .C(N9211), .D(n3670), .Z(
        n2402) );
  CND3XL U10427 ( .A(n2405), .B(n2406), .C(n2407), .Z(N10254) );
  CANR2X1 U10428 ( .A(N3006), .B(n3600), .C(n3634), .D(N7349), .Z(n2407) );
  CND2X1 U10429 ( .A(N6088), .B(n3698), .Z(n2406) );
  CANR2X1 U10430 ( .A(mem_data1[930]), .B(n3898), .C(N9210), .D(n3670), .Z(
        n2405) );
  CND3XL U10431 ( .A(n2408), .B(n2409), .C(n2410), .Z(N10253) );
  CND3XL U10432 ( .A(n2411), .B(n2412), .C(n2413), .Z(N10252) );
  CANR2X1 U10433 ( .A(N3004), .B(n3600), .C(n3634), .D(N7351), .Z(n2413) );
  CND2X1 U10434 ( .A(N6086), .B(n3685), .Z(n2412) );
  CANR2X1 U10435 ( .A(mem_data1[928]), .B(n3898), .C(N9208), .D(n3670), .Z(
        n2411) );
  CND3XL U10436 ( .A(n2414), .B(n2415), .C(n2416), .Z(N10251) );
  CANR2X1 U10437 ( .A(N3003), .B(n3600), .C(n3634), .D(N7352), .Z(n2416) );
  CND2X1 U10438 ( .A(N6085), .B(n3696), .Z(n2415) );
  CANR2X1 U10439 ( .A(mem_data1[927]), .B(n3898), .C(N9207), .D(n3670), .Z(
        n2414) );
  CND3XL U10440 ( .A(n2417), .B(n2418), .C(n2419), .Z(N10250) );
  CANR2X1 U10441 ( .A(N3002), .B(n3600), .C(n3634), .D(N7353), .Z(n2419) );
  CND2X1 U10442 ( .A(N6084), .B(n3698), .Z(n2418) );
  CANR2X1 U10443 ( .A(mem_data1[926]), .B(n3898), .C(N9206), .D(n3670), .Z(
        n2417) );
  CND3XL U10444 ( .A(n2420), .B(n2421), .C(n2422), .Z(N10249) );
  CANR2X1 U10445 ( .A(N3001), .B(n3600), .C(n3634), .D(N7354), .Z(n2422) );
  CND2X1 U10446 ( .A(N6083), .B(n3684), .Z(n2421) );
  CANR2X1 U10447 ( .A(mem_data1[925]), .B(n3898), .C(N9205), .D(n3670), .Z(
        n2420) );
  CND3XL U10448 ( .A(n2423), .B(n2424), .C(n2425), .Z(N10248) );
  CANR2X1 U10449 ( .A(N3000), .B(n3600), .C(n3634), .D(N7355), .Z(n2425) );
  CND2X1 U10450 ( .A(N6082), .B(n3695), .Z(n2424) );
  CANR2X1 U10451 ( .A(mem_data1[924]), .B(n3898), .C(N9204), .D(n3670), .Z(
        n2423) );
  CND3XL U10452 ( .A(n2426), .B(n2427), .C(n2428), .Z(N10247) );
  CANR2X1 U10453 ( .A(N2999), .B(n3600), .C(n3634), .D(N7356), .Z(n2428) );
  CND2X1 U10454 ( .A(N6081), .B(n3690), .Z(n2427) );
  CANR2X1 U10455 ( .A(mem_data1[923]), .B(n3898), .C(N9203), .D(n3670), .Z(
        n2426) );
  CND3XL U10456 ( .A(n2429), .B(n2430), .C(n2431), .Z(N10246) );
  CANR2X1 U10457 ( .A(N2998), .B(n3600), .C(n3634), .D(N7357), .Z(n2431) );
  CND2X1 U10458 ( .A(N6080), .B(n3692), .Z(n2430) );
  CANR2X1 U10459 ( .A(mem_data1[922]), .B(n3898), .C(N9202), .D(n3670), .Z(
        n2429) );
  CND3XL U10460 ( .A(n2432), .B(n2433), .C(n2434), .Z(N10245) );
  CANR2X1 U10461 ( .A(N2997), .B(n3600), .C(n3634), .D(N7358), .Z(n2434) );
  CND2X1 U10462 ( .A(N6079), .B(n3687), .Z(n2433) );
  CANR2X1 U10463 ( .A(mem_data1[921]), .B(n3898), .C(N9201), .D(n3670), .Z(
        n2432) );
  CND3XL U10464 ( .A(n2435), .B(n2436), .C(n2437), .Z(N10244) );
  CANR2X1 U10465 ( .A(N2996), .B(n3600), .C(n3634), .D(N7359), .Z(n2437) );
  CND2X1 U10466 ( .A(N6078), .B(n3686), .Z(n2436) );
  CANR2X1 U10467 ( .A(mem_data1[920]), .B(n3898), .C(N9200), .D(n3670), .Z(
        n2435) );
  CND3XL U10468 ( .A(n2438), .B(n2439), .C(n2440), .Z(N10243) );
  CANR2X1 U10469 ( .A(N2995), .B(n3600), .C(n3633), .D(N7360), .Z(n2440) );
  CND2X1 U10470 ( .A(N6077), .B(n3693), .Z(n2439) );
  CANR2X1 U10471 ( .A(mem_data1[919]), .B(n3898), .C(N9199), .D(n3670), .Z(
        n2438) );
  CND3XL U10472 ( .A(n2441), .B(n2442), .C(n2443), .Z(N10242) );
  CANR2X1 U10473 ( .A(N2994), .B(n3600), .C(n3633), .D(N7361), .Z(n2443) );
  CND2X1 U10474 ( .A(N6076), .B(n3683), .Z(n2442) );
  CANR2X1 U10475 ( .A(mem_data1[918]), .B(n3898), .C(N9198), .D(n3670), .Z(
        n2441) );
  CND3XL U10476 ( .A(n2444), .B(n2445), .C(n2446), .Z(N10241) );
  CANR2X1 U10477 ( .A(N2993), .B(n3600), .C(n3633), .D(N7362), .Z(n2446) );
  CND2X1 U10478 ( .A(N6075), .B(n3685), .Z(n2445) );
  CANR2X1 U10479 ( .A(mem_data1[917]), .B(n3898), .C(N9197), .D(n3670), .Z(
        n2444) );
  CND3XL U10480 ( .A(n2447), .B(n2448), .C(n2449), .Z(N10240) );
  CANR2X1 U10481 ( .A(N2992), .B(n3600), .C(n3633), .D(N7363), .Z(n2449) );
  CND2X1 U10482 ( .A(N6074), .B(n3697), .Z(n2448) );
  CANR2X1 U10483 ( .A(mem_data1[916]), .B(n3898), .C(N9196), .D(n3671), .Z(
        n2447) );
  CND3XL U10484 ( .A(n2450), .B(n2451), .C(n2452), .Z(N10239) );
  CANR2X1 U10485 ( .A(N2991), .B(n3600), .C(n3633), .D(N7364), .Z(n2452) );
  CND2X1 U10486 ( .A(N6073), .B(n3698), .Z(n2451) );
  CANR2X1 U10487 ( .A(mem_data1[915]), .B(n3898), .C(N9195), .D(n3676), .Z(
        n2450) );
  CND3XL U10488 ( .A(n2453), .B(n2454), .C(n2455), .Z(N10238) );
  CND3XL U10489 ( .A(n2456), .B(n2457), .C(n2458), .Z(N10237) );
  CND2X1 U10490 ( .A(N6071), .B(n3691), .Z(n2457) );
  CND3XL U10491 ( .A(n2459), .B(n2460), .C(n2461), .Z(N10236) );
  CANR2X1 U10492 ( .A(N2988), .B(n3599), .C(n3633), .D(N7367), .Z(n2461) );
  CND2X1 U10493 ( .A(N6070), .B(n3690), .Z(n2460) );
  CND3XL U10494 ( .A(n2462), .B(n2463), .C(n2464), .Z(N10235) );
  CND2X1 U10495 ( .A(N6069), .B(n3690), .Z(n2463) );
  CND3XL U10496 ( .A(n2465), .B(n2466), .C(n2467), .Z(N10234) );
  CND2X1 U10497 ( .A(N6068), .B(n3696), .Z(n2466) );
  CND3XL U10498 ( .A(n2468), .B(n2469), .C(n2470), .Z(N10233) );
  CND2X1 U10499 ( .A(N6067), .B(n3694), .Z(n2469) );
  CND3XL U10500 ( .A(n2471), .B(n2472), .C(n2473), .Z(N10232) );
  CND2X1 U10501 ( .A(N6066), .B(n3695), .Z(n2472) );
  CND3XL U10502 ( .A(n2474), .B(n2475), .C(n2476), .Z(N10231) );
  CND2X1 U10503 ( .A(N6065), .B(n3697), .Z(n2475) );
  CND3XL U10504 ( .A(n2477), .B(n2478), .C(n2479), .Z(N10230) );
  CND3XL U10505 ( .A(n2480), .B(n2481), .C(n2482), .Z(N10229) );
  CND3XL U10506 ( .A(n2483), .B(n2484), .C(n2485), .Z(N10228) );
  CND3XL U10507 ( .A(n2486), .B(n2487), .C(n2488), .Z(N10227) );
  CND3XL U10508 ( .A(n2489), .B(n2490), .C(n2491), .Z(N10226) );
  CANR2X1 U10509 ( .A(N2978), .B(n3601), .C(n3635), .D(N7377), .Z(n2491) );
  CND2X1 U10510 ( .A(N6060), .B(n3684), .Z(n2490) );
  CANR2X1 U10511 ( .A(mem_data1[902]), .B(n3898), .C(N9182), .D(n3673), .Z(
        n2489) );
  CND3XL U10512 ( .A(n2492), .B(n2493), .C(n2494), .Z(N10225) );
  CANR2X1 U10513 ( .A(N2977), .B(n3601), .C(n3635), .D(N7378), .Z(n2494) );
  CND2X1 U10514 ( .A(N6059), .B(n3695), .Z(n2493) );
  CANR2X1 U10515 ( .A(mem_data1[901]), .B(n3898), .C(N9181), .D(n3673), .Z(
        n2492) );
  CND3XL U10516 ( .A(n2495), .B(n2496), .C(n2497), .Z(N10224) );
  CANR2X1 U10517 ( .A(N2976), .B(n3601), .C(n3635), .D(N7379), .Z(n2497) );
  CND2X1 U10518 ( .A(N6058), .B(n3687), .Z(n2496) );
  CANR2X1 U10519 ( .A(mem_data1[900]), .B(n3898), .C(N9180), .D(n3673), .Z(
        n2495) );
  CND3XL U10520 ( .A(n2498), .B(n2499), .C(n2500), .Z(N10223) );
  CANR2X1 U10521 ( .A(N2975), .B(n3601), .C(n3635), .D(N7380), .Z(n2500) );
  CND2X1 U10522 ( .A(N6057), .B(n3695), .Z(n2499) );
  CANR2X1 U10523 ( .A(mem_data1[899]), .B(n3898), .C(N9179), .D(n3673), .Z(
        n2498) );
  CND3XL U10524 ( .A(n2501), .B(n2502), .C(n2503), .Z(N10222) );
  CANR2X1 U10525 ( .A(N2974), .B(n3601), .C(n3635), .D(N7381), .Z(n2503) );
  CND2X1 U10526 ( .A(N6056), .B(n3686), .Z(n2502) );
  CANR2X1 U10527 ( .A(mem_data1[898]), .B(n3898), .C(N9178), .D(n3673), .Z(
        n2501) );
  CND3XL U10528 ( .A(n2504), .B(n2505), .C(n2506), .Z(N10221) );
  CANR2X1 U10529 ( .A(N2973), .B(n3601), .C(n3635), .D(N7382), .Z(n2506) );
  CND2X1 U10530 ( .A(N6055), .B(n3693), .Z(n2505) );
  CANR2X1 U10531 ( .A(mem_data1[897]), .B(n3898), .C(N9177), .D(n3673), .Z(
        n2504) );
  CND3XL U10532 ( .A(n2507), .B(n2508), .C(n2509), .Z(N10220) );
  CANR2X1 U10533 ( .A(N2972), .B(n3601), .C(n3635), .D(N7383), .Z(n2509) );
  CND2X1 U10534 ( .A(N6054), .B(n3698), .Z(n2508) );
  CANR2X1 U10535 ( .A(mem_data1[896]), .B(n3898), .C(N9176), .D(n3672), .Z(
        n2507) );
  CND3XL U10536 ( .A(n2510), .B(n2511), .C(n2512), .Z(N10219) );
  CANR2X1 U10537 ( .A(N2971), .B(n3601), .C(n3635), .D(N7384), .Z(n2512) );
  CND2X1 U10538 ( .A(N6053), .B(n3687), .Z(n2511) );
  CANR2X1 U10539 ( .A(mem_data1[895]), .B(n3898), .C(N9175), .D(n3672), .Z(
        n2510) );
  CND3XL U10540 ( .A(n2513), .B(n2514), .C(n2515), .Z(N10218) );
  CANR2X1 U10541 ( .A(N2970), .B(n3601), .C(n3635), .D(N7385), .Z(n2515) );
  CND2X1 U10542 ( .A(N6052), .B(n3697), .Z(n2514) );
  CANR2X1 U10543 ( .A(mem_data1[894]), .B(n3898), .C(N9174), .D(n3670), .Z(
        n2513) );
  CND3XL U10544 ( .A(n2516), .B(n2517), .C(n2518), .Z(N10217) );
  CANR2X1 U10545 ( .A(N2969), .B(n3601), .C(n3635), .D(N7386), .Z(n2518) );
  CND2X1 U10546 ( .A(N6051), .B(n3694), .Z(n2517) );
  CANR2X1 U10547 ( .A(mem_data1[893]), .B(n3898), .C(N9173), .D(n3663), .Z(
        n2516) );
  CND3XL U10548 ( .A(n2519), .B(n2520), .C(n2521), .Z(N10216) );
  CANR2X1 U10549 ( .A(N2968), .B(n3601), .C(n3634), .D(N7387), .Z(n2521) );
  CND2X1 U10550 ( .A(N6050), .B(n3691), .Z(n2520) );
  CANR2X1 U10551 ( .A(mem_data1[892]), .B(n3898), .C(N9172), .D(n3663), .Z(
        n2519) );
  CND3XL U10552 ( .A(n2522), .B(n2523), .C(n2524), .Z(N10215) );
  CANR2X1 U10553 ( .A(N2967), .B(n3601), .C(n3634), .D(N7388), .Z(n2524) );
  CND2X1 U10554 ( .A(N6049), .B(n3694), .Z(n2523) );
  CANR2X1 U10555 ( .A(mem_data1[891]), .B(n3898), .C(N9171), .D(n3664), .Z(
        n2522) );
  CND3XL U10556 ( .A(n2525), .B(n2526), .C(n2527), .Z(N10214) );
  CANR2X1 U10557 ( .A(N2966), .B(n3601), .C(n3634), .D(N7389), .Z(n2527) );
  CND2X1 U10558 ( .A(N6048), .B(n3683), .Z(n2526) );
  CANR2X1 U10559 ( .A(mem_data1[890]), .B(n3898), .C(N9170), .D(n3664), .Z(
        n2525) );
  CND3XL U10560 ( .A(n2528), .B(n2529), .C(n2530), .Z(N10213) );
  CANR2X1 U10561 ( .A(N2965), .B(n3601), .C(n3634), .D(N7390), .Z(n2530) );
  CND2X1 U10562 ( .A(N6047), .B(n3696), .Z(n2529) );
  CANR2X1 U10563 ( .A(mem_data1[889]), .B(n3898), .C(N9169), .D(n3664), .Z(
        n2528) );
  CND3XL U10564 ( .A(n2531), .B(n2532), .C(n2533), .Z(N10212) );
  CANR2X1 U10565 ( .A(N2964), .B(n3601), .C(n3634), .D(N7391), .Z(n2533) );
  CND2X1 U10566 ( .A(N6046), .B(n3695), .Z(n2532) );
  CANR2X1 U10567 ( .A(mem_data1[888]), .B(n3898), .C(N9168), .D(n3664), .Z(
        n2531) );
  CND3XL U10568 ( .A(n2534), .B(n2535), .C(n2536), .Z(N10211) );
  CANR2X1 U10569 ( .A(N2963), .B(n3600), .C(n3634), .D(N7392), .Z(n2536) );
  CND2X1 U10570 ( .A(N6045), .B(n3690), .Z(n2535) );
  CANR2X1 U10571 ( .A(mem_data1[887]), .B(n3898), .C(N9167), .D(n3664), .Z(
        n2534) );
  CND3XL U10572 ( .A(n2537), .B(n2538), .C(n2539), .Z(N10210) );
  CANR2X1 U10573 ( .A(N2962), .B(n3600), .C(n3634), .D(N7393), .Z(n2539) );
  CND2X1 U10574 ( .A(N6044), .B(n3694), .Z(n2538) );
  CANR2X1 U10575 ( .A(mem_data1[886]), .B(n3898), .C(N9166), .D(n3664), .Z(
        n2537) );
  CND3XL U10576 ( .A(n2540), .B(n2541), .C(n2542), .Z(N10209) );
  CANR2X1 U10577 ( .A(N2961), .B(n3575), .C(n3634), .D(N7394), .Z(n2542) );
  CND2X1 U10578 ( .A(N6043), .B(n3691), .Z(n2541) );
  CANR2X1 U10579 ( .A(mem_data1[885]), .B(n3898), .C(N9165), .D(n3664), .Z(
        n2540) );
  CND3XL U10580 ( .A(n2543), .B(n2544), .C(n2545), .Z(N10208) );
  CANR2X1 U10581 ( .A(N2960), .B(n3575), .C(n3634), .D(N7395), .Z(n2545) );
  CND2X1 U10582 ( .A(N6042), .B(n3695), .Z(n2544) );
  CANR2X1 U10583 ( .A(mem_data1[884]), .B(n3898), .C(N9164), .D(n3664), .Z(
        n2543) );
  CND3XL U10584 ( .A(n2546), .B(n2547), .C(n2548), .Z(N10207) );
  CANR2X1 U10585 ( .A(N2959), .B(n3575), .C(n3634), .D(N7396), .Z(n2548) );
  CND2X1 U10586 ( .A(N6041), .B(n3684), .Z(n2547) );
  CANR2X1 U10587 ( .A(mem_data1[883]), .B(n3898), .C(N9163), .D(n3664), .Z(
        n2546) );
  CND3XL U10588 ( .A(n2549), .B(n2550), .C(n2551), .Z(N10206) );
  CANR2X1 U10589 ( .A(N2958), .B(n3575), .C(n3634), .D(N7397), .Z(n2551) );
  CND2X1 U10590 ( .A(N6040), .B(n3684), .Z(n2550) );
  CANR2X1 U10591 ( .A(mem_data1[882]), .B(n3898), .C(N9162), .D(n3664), .Z(
        n2549) );
  CND3XL U10592 ( .A(n2552), .B(n2553), .C(n2554), .Z(N10205) );
  CANR2X1 U10593 ( .A(N2957), .B(n3575), .C(n3634), .D(N7398), .Z(n2554) );
  CND2X1 U10594 ( .A(N6039), .B(n3686), .Z(n2553) );
  CANR2X1 U10595 ( .A(mem_data1[881]), .B(n3898), .C(N9161), .D(n3664), .Z(
        n2552) );
  CND3XL U10596 ( .A(n2555), .B(n2556), .C(n2557), .Z(N10204) );
  CANR2X1 U10597 ( .A(N2956), .B(n3575), .C(n3634), .D(N7399), .Z(n2557) );
  CND2X1 U10598 ( .A(N6038), .B(n3687), .Z(n2556) );
  CANR2X1 U10599 ( .A(mem_data1[880]), .B(n3898), .C(N9160), .D(n3664), .Z(
        n2555) );
  CND3XL U10600 ( .A(n2558), .B(n2559), .C(n2560), .Z(N10203) );
  CANR2X1 U10601 ( .A(N2955), .B(n3575), .C(n3611), .D(N7400), .Z(n2560) );
  CND2X1 U10602 ( .A(N6037), .B(n3694), .Z(n2559) );
  CANR2X1 U10603 ( .A(mem_data1[879]), .B(n3898), .C(N9159), .D(n3664), .Z(
        n2558) );
  CND3XL U10604 ( .A(n2561), .B(n2562), .C(n2563), .Z(N10202) );
  CANR2X1 U10605 ( .A(N2954), .B(n3574), .C(n3611), .D(N7401), .Z(n2563) );
  CND2X1 U10606 ( .A(N6036), .B(n3689), .Z(n2562) );
  CANR2X1 U10607 ( .A(mem_data1[878]), .B(n3898), .C(N9158), .D(n3664), .Z(
        n2561) );
  CND3XL U10608 ( .A(n2564), .B(n2565), .C(n2566), .Z(N10201) );
  CANR2X1 U10609 ( .A(N2953), .B(n3574), .C(n3611), .D(N7402), .Z(n2566) );
  CND2X1 U10610 ( .A(N6035), .B(n3694), .Z(n2565) );
  CANR2X1 U10611 ( .A(mem_data1[877]), .B(n3898), .C(N9157), .D(n3664), .Z(
        n2564) );
  CND3XL U10612 ( .A(n2567), .B(n2568), .C(n2569), .Z(N10200) );
  CANR2X1 U10613 ( .A(N2952), .B(n3574), .C(n3611), .D(N7403), .Z(n2569) );
  CND2X1 U10614 ( .A(N6034), .B(n3690), .Z(n2568) );
  CANR2X1 U10615 ( .A(mem_data1[876]), .B(n3898), .C(N9156), .D(n3664), .Z(
        n2567) );
  CND3XL U10616 ( .A(n2570), .B(n2571), .C(n2572), .Z(N10199) );
  CANR2X1 U10617 ( .A(N2951), .B(n3574), .C(n3611), .D(N7404), .Z(n2572) );
  CND2X1 U10618 ( .A(N6033), .B(n3690), .Z(n2571) );
  CANR2X1 U10619 ( .A(mem_data1[875]), .B(n3898), .C(N9155), .D(n3664), .Z(
        n2570) );
  CND3XL U10620 ( .A(n2573), .B(n2574), .C(n2575), .Z(N10198) );
  CANR2X1 U10621 ( .A(N2950), .B(n3574), .C(n3610), .D(N7405), .Z(n2575) );
  CND2X1 U10622 ( .A(N6032), .B(n3697), .Z(n2574) );
  CANR2X1 U10623 ( .A(mem_data1[874]), .B(n3898), .C(N9154), .D(n3664), .Z(
        n2573) );
  CND3XL U10624 ( .A(n2576), .B(n2577), .C(n2578), .Z(N10197) );
  CND3XL U10625 ( .A(n2579), .B(n2580), .C(n2581), .Z(N10196) );
  CND3XL U10626 ( .A(n2582), .B(n2583), .C(n2584), .Z(N10195) );
  CANR2X1 U10627 ( .A(N2947), .B(n3574), .C(n3610), .D(N7408), .Z(n2584) );
  CND2X1 U10628 ( .A(N6029), .B(n3689), .Z(n2583) );
  CANR2X1 U10629 ( .A(mem_data1[871]), .B(n3898), .C(N9151), .D(n3662), .Z(
        n2582) );
  CND3XL U10630 ( .A(n2585), .B(n2586), .C(n2587), .Z(N10194) );
  CANR2X1 U10631 ( .A(N2946), .B(n3574), .C(n3610), .D(N7409), .Z(n2587) );
  CND2X1 U10632 ( .A(N6028), .B(n3693), .Z(n2586) );
  CANR2X1 U10633 ( .A(mem_data1[870]), .B(n3898), .C(N9150), .D(n3662), .Z(
        n2585) );
  CND3XL U10634 ( .A(n2588), .B(n2589), .C(n2590), .Z(N10193) );
  CANR2X1 U10635 ( .A(N2945), .B(n3574), .C(n3610), .D(N7410), .Z(n2590) );
  CND2X1 U10636 ( .A(N6027), .B(n3684), .Z(n2589) );
  CANR2X1 U10637 ( .A(mem_data1[869]), .B(n3898), .C(N9149), .D(n3663), .Z(
        n2588) );
  CND3XL U10638 ( .A(n2591), .B(n2592), .C(n2593), .Z(N10192) );
  CANR2X1 U10639 ( .A(N2944), .B(n3574), .C(n3610), .D(N7411), .Z(n2593) );
  CND2X1 U10640 ( .A(N6026), .B(n3685), .Z(n2592) );
  CANR2X1 U10641 ( .A(mem_data1[868]), .B(n3898), .C(N9148), .D(n3663), .Z(
        n2591) );
  CND3XL U10642 ( .A(n2594), .B(n2595), .C(n2596), .Z(N10191) );
  CANR2X1 U10643 ( .A(N2943), .B(n3574), .C(n3610), .D(N7412), .Z(n2596) );
  CND2X1 U10644 ( .A(N6025), .B(n3695), .Z(n2595) );
  CANR2X1 U10645 ( .A(mem_data1[867]), .B(n3898), .C(N9147), .D(n3663), .Z(
        n2594) );
  CND3XL U10646 ( .A(n2597), .B(n2598), .C(n2599), .Z(N10190) );
  CANR2X1 U10647 ( .A(N2942), .B(n3576), .C(n3610), .D(N7413), .Z(n2599) );
  CND2X1 U10648 ( .A(N6024), .B(n3688), .Z(n2598) );
  CANR2X1 U10649 ( .A(mem_data1[866]), .B(n3898), .C(N9146), .D(n3663), .Z(
        n2597) );
  CND3XL U10650 ( .A(n2600), .B(n2601), .C(n2602), .Z(N10189) );
  CANR2X1 U10651 ( .A(N2941), .B(n3578), .C(n3610), .D(N7414), .Z(n2602) );
  CND2X1 U10652 ( .A(N6023), .B(n3686), .Z(n2601) );
  CANR2X1 U10653 ( .A(mem_data1[865]), .B(n3898), .C(N9145), .D(n3663), .Z(
        n2600) );
  CND3XL U10654 ( .A(n2603), .B(n2604), .C(n2605), .Z(N10188) );
  CANR2X1 U10655 ( .A(N2940), .B(n3597), .C(n3610), .D(N7415), .Z(n2605) );
  CND2X1 U10656 ( .A(N6022), .B(n3698), .Z(n2604) );
  CANR2X1 U10657 ( .A(mem_data1[864]), .B(n3898), .C(N9144), .D(n3663), .Z(
        n2603) );
  CND3XL U10658 ( .A(n2606), .B(n2607), .C(n2608), .Z(N10187) );
  CANR2X1 U10659 ( .A(N2939), .B(n3601), .C(n3610), .D(N7416), .Z(n2608) );
  CND2X1 U10660 ( .A(N6021), .B(n3697), .Z(n2607) );
  CANR2X1 U10661 ( .A(mem_data1[863]), .B(n3898), .C(N9143), .D(n3663), .Z(
        n2606) );
  CND3XL U10662 ( .A(n2609), .B(n2610), .C(n2611), .Z(N10186) );
  CANR2X1 U10663 ( .A(N2938), .B(n3601), .C(n3610), .D(N7417), .Z(n2611) );
  CND2X1 U10664 ( .A(N6020), .B(n3687), .Z(n2610) );
  CANR2X1 U10665 ( .A(mem_data1[862]), .B(n3898), .C(N9142), .D(n3663), .Z(
        n2609) );
  CND3XL U10666 ( .A(n2612), .B(n2613), .C(n2614), .Z(N10185) );
  CANR2X1 U10667 ( .A(N2937), .B(n3576), .C(n3610), .D(N7418), .Z(n2614) );
  CND2X1 U10668 ( .A(N6019), .B(n3684), .Z(n2613) );
  CANR2X1 U10669 ( .A(mem_data1[861]), .B(n3898), .C(N9141), .D(n3663), .Z(
        n2612) );
  CND3XL U10670 ( .A(n2615), .B(n2616), .C(n2617), .Z(N10184) );
  CANR2X1 U10671 ( .A(N2936), .B(n3576), .C(n3610), .D(N7419), .Z(n2617) );
  CND2X1 U10672 ( .A(N6018), .B(n3696), .Z(n2616) );
  CANR2X1 U10673 ( .A(mem_data1[860]), .B(n3898), .C(N9140), .D(n3663), .Z(
        n2615) );
  CND3XL U10674 ( .A(n2618), .B(n2619), .C(n2620), .Z(N10183) );
  CANR2X1 U10675 ( .A(N2935), .B(n3576), .C(n3610), .D(N7420), .Z(n2620) );
  CND2X1 U10676 ( .A(N6017), .B(n3695), .Z(n2619) );
  CANR2X1 U10677 ( .A(mem_data1[859]), .B(n3898), .C(N9139), .D(n3663), .Z(
        n2618) );
  CND3XL U10678 ( .A(n2621), .B(n2622), .C(n2623), .Z(N10182) );
  CANR2X1 U10679 ( .A(N2934), .B(n3576), .C(n3610), .D(N7421), .Z(n2623) );
  CND2X1 U10680 ( .A(N6016), .B(n3690), .Z(n2622) );
  CANR2X1 U10681 ( .A(mem_data1[858]), .B(n3898), .C(N9138), .D(n3663), .Z(
        n2621) );
  CND3XL U10682 ( .A(n2624), .B(n2625), .C(n2626), .Z(N10181) );
  CANR2X1 U10683 ( .A(N2933), .B(n3576), .C(n3610), .D(N7422), .Z(n2626) );
  CND2X1 U10684 ( .A(N6015), .B(n3694), .Z(n2625) );
  CANR2X1 U10685 ( .A(mem_data1[857]), .B(n3898), .C(N9137), .D(n3663), .Z(
        n2624) );
  CND3XL U10686 ( .A(n2627), .B(n2628), .C(n2629), .Z(N10180) );
  CANR2X1 U10687 ( .A(N2932), .B(n3576), .C(n3610), .D(N7423), .Z(n2629) );
  CND2X1 U10688 ( .A(N6014), .B(n3691), .Z(n2628) );
  CANR2X1 U10689 ( .A(mem_data1[856]), .B(n3898), .C(N9136), .D(n3663), .Z(
        n2627) );
  CND3XL U10690 ( .A(n2630), .B(n2631), .C(n2632), .Z(N10179) );
  CANR2X1 U10691 ( .A(N2931), .B(n3576), .C(n3610), .D(N7424), .Z(n2632) );
  CND2X1 U10692 ( .A(N6013), .B(n3698), .Z(n2631) );
  CANR2X1 U10693 ( .A(mem_data1[855]), .B(n3898), .C(N9135), .D(n3663), .Z(
        n2630) );
  CND3XL U10694 ( .A(n2633), .B(n2634), .C(n2635), .Z(N10178) );
  CANR2X1 U10695 ( .A(N2930), .B(n3575), .C(n3610), .D(N7425), .Z(n2635) );
  CND2X1 U10696 ( .A(N6012), .B(n3691), .Z(n2634) );
  CANR2X1 U10697 ( .A(mem_data1[854]), .B(n3898), .C(N9134), .D(n3663), .Z(
        n2633) );
  CND3XL U10698 ( .A(n2636), .B(n2637), .C(n2638), .Z(N10177) );
  CANR2X1 U10699 ( .A(N2929), .B(n3575), .C(n3612), .D(N7426), .Z(n2638) );
  CND2X1 U10700 ( .A(N6011), .B(n3696), .Z(n2637) );
  CANR2X1 U10701 ( .A(mem_data1[853]), .B(n3898), .C(N9133), .D(n3663), .Z(
        n2636) );
  CND3XL U10702 ( .A(n2639), .B(n2640), .C(n2641), .Z(N10176) );
  CANR2X1 U10703 ( .A(N2928), .B(n3575), .C(n3612), .D(N7427), .Z(n2641) );
  CND2X1 U10704 ( .A(N6010), .B(n3695), .Z(n2640) );
  CANR2X1 U10705 ( .A(mem_data1[852]), .B(n3898), .C(N9132), .D(n3663), .Z(
        n2639) );
  CND3XL U10706 ( .A(n2642), .B(n2643), .C(n2644), .Z(N10175) );
  CANR2X1 U10707 ( .A(N2927), .B(n3575), .C(n3612), .D(N7428), .Z(n2644) );
  CND2X1 U10708 ( .A(N6009), .B(n3690), .Z(n2643) );
  CANR2X1 U10709 ( .A(mem_data1[851]), .B(n3898), .C(N9131), .D(n3663), .Z(
        n2642) );
  CND3XL U10710 ( .A(n2645), .B(n2646), .C(n2647), .Z(N10174) );
  CANR2X1 U10711 ( .A(N2926), .B(n3575), .C(n3612), .D(N7429), .Z(n2647) );
  CND2X1 U10712 ( .A(N6008), .B(n3694), .Z(n2646) );
  CANR2X1 U10713 ( .A(mem_data1[850]), .B(n3898), .C(N9130), .D(n3663), .Z(
        n2645) );
  CND3XL U10714 ( .A(n2648), .B(n2649), .C(n2650), .Z(N10173) );
  CND3XL U10715 ( .A(n2651), .B(n2652), .C(n2653), .Z(N10172) );
  CANR2X1 U10716 ( .A(N2924), .B(n3575), .C(n3611), .D(N7431), .Z(n2653) );
  CND3XL U10717 ( .A(n2654), .B(n2655), .C(n2656), .Z(N10171) );
  CND3XL U10718 ( .A(n2657), .B(n2658), .C(n2659), .Z(N10170) );
  CND3XL U10719 ( .A(n2660), .B(n2661), .C(n2662), .Z(N10169) );
  CND3XL U10720 ( .A(n2663), .B(n2664), .C(n2665), .Z(N10168) );
  CND3XL U10721 ( .A(n2666), .B(n2667), .C(n2668), .Z(N10167) );
  CND3XL U10722 ( .A(n2669), .B(n2670), .C(n2671), .Z(N10166) );
  CND3XL U10723 ( .A(n2672), .B(n2673), .C(n2674), .Z(N10165) );
  CND3XL U10724 ( .A(n2675), .B(n2676), .C(n2677), .Z(N10164) );
  CND3XL U10725 ( .A(n2678), .B(n2679), .C(n2680), .Z(N10163) );
  CND3XL U10726 ( .A(n2681), .B(n2682), .C(n2683), .Z(N10162) );
  CND3XL U10727 ( .A(n2684), .B(n2685), .C(n2686), .Z(N10161) );
  CND3XL U10728 ( .A(n2687), .B(n2688), .C(n2689), .Z(N10160) );
  CND3XL U10729 ( .A(n2690), .B(n2691), .C(n2692), .Z(N10159) );
  CND3XL U10730 ( .A(n2693), .B(n2694), .C(n2695), .Z(N10158) );
  CND3XL U10731 ( .A(n2696), .B(n2697), .C(n2698), .Z(N10157) );
  CND3XL U10732 ( .A(n2699), .B(n2700), .C(n2701), .Z(N10156) );
  CANR2X1 U10733 ( .A(N2908), .B(n3577), .C(n3611), .D(N7447), .Z(n2701) );
  CND2X1 U10734 ( .A(N5990), .B(n3689), .Z(n2700) );
  CANR2X1 U10735 ( .A(mem_data1[832]), .B(n3898), .C(N9112), .D(n3662), .Z(
        n2699) );
  CND3XL U10736 ( .A(n2702), .B(n2703), .C(n2704), .Z(N10155) );
  CANR2X1 U10737 ( .A(N2907), .B(n3577), .C(n3611), .D(N7448), .Z(n2704) );
  CND2X1 U10738 ( .A(N5989), .B(n3694), .Z(n2703) );
  CANR2X1 U10739 ( .A(mem_data1[831]), .B(n3898), .C(N9111), .D(n3662), .Z(
        n2702) );
  CND3XL U10740 ( .A(n2705), .B(n2706), .C(n2707), .Z(N10154) );
  CANR2X1 U10741 ( .A(N2906), .B(n3577), .C(n3611), .D(N7449), .Z(n2707) );
  CND2X1 U10742 ( .A(N5988), .B(n3696), .Z(n2706) );
  CANR2X1 U10743 ( .A(mem_data1[830]), .B(n3898), .C(N9110), .D(n3662), .Z(
        n2705) );
  CND3XL U10744 ( .A(n2708), .B(n2709), .C(n2710), .Z(N10153) );
  CANR2X1 U10745 ( .A(N2905), .B(n3577), .C(n3611), .D(N7450), .Z(n2710) );
  CND2X1 U10746 ( .A(N5987), .B(n3683), .Z(n2709) );
  CANR2X1 U10747 ( .A(mem_data1[829]), .B(n3898), .C(N9109), .D(n3662), .Z(
        n2708) );
  CND3XL U10748 ( .A(n2711), .B(n2712), .C(n2713), .Z(N10152) );
  CANR2X1 U10749 ( .A(N2904), .B(n3576), .C(n3611), .D(N7451), .Z(n2713) );
  CND2X1 U10750 ( .A(N5986), .B(n3691), .Z(n2712) );
  CANR2X1 U10751 ( .A(mem_data1[828]), .B(n3898), .C(N9108), .D(n3662), .Z(
        n2711) );
  CND3XL U10752 ( .A(n2714), .B(n2715), .C(n2716), .Z(N10151) );
  CANR2X1 U10753 ( .A(N2903), .B(n3576), .C(n3611), .D(N7452), .Z(n2716) );
  CND2X1 U10754 ( .A(N5985), .B(n3685), .Z(n2715) );
  CANR2X1 U10755 ( .A(mem_data1[827]), .B(n3898), .C(N9107), .D(n3660), .Z(
        n2714) );
  CND3XL U10756 ( .A(n2717), .B(n2718), .C(n2719), .Z(N10150) );
  CANR2X1 U10757 ( .A(N2902), .B(n3576), .C(n3613), .D(N7453), .Z(n2719) );
  CND2X1 U10758 ( .A(N5984), .B(n3697), .Z(n2718) );
  CANR2X1 U10759 ( .A(mem_data1[826]), .B(n3898), .C(N9106), .D(n3660), .Z(
        n2717) );
  CND3XL U10760 ( .A(n2720), .B(n2721), .C(n2722), .Z(N10149) );
  CANR2X1 U10761 ( .A(N2901), .B(n3576), .C(n3613), .D(N7454), .Z(n2722) );
  CND2X1 U10762 ( .A(N5983), .B(n3698), .Z(n2721) );
  CANR2X1 U10763 ( .A(mem_data1[825]), .B(n3898), .C(N9105), .D(n3660), .Z(
        n2720) );
  CND3XL U10764 ( .A(n2723), .B(n2724), .C(n2725), .Z(N10148) );
  CANR2X1 U10765 ( .A(N2900), .B(n3576), .C(n3613), .D(N7455), .Z(n2725) );
  CND2X1 U10766 ( .A(N5982), .B(n3689), .Z(n2724) );
  CANR2X1 U10767 ( .A(mem_data1[824]), .B(n3898), .C(N9104), .D(n3661), .Z(
        n2723) );
  CND3XL U10768 ( .A(n2726), .B(n2727), .C(n2728), .Z(N10147) );
  CANR2X1 U10769 ( .A(N2899), .B(n3576), .C(n3613), .D(N7456), .Z(n2728) );
  CND2X1 U10770 ( .A(N5981), .B(n3688), .Z(n2727) );
  CANR2X1 U10771 ( .A(mem_data1[823]), .B(n3898), .C(N9103), .D(n3661), .Z(
        n2726) );
  CND3XL U10772 ( .A(n2729), .B(n2730), .C(n2731), .Z(N10146) );
  CANR2X1 U10773 ( .A(N2898), .B(n3576), .C(n3613), .D(N7457), .Z(n2731) );
  CND2X1 U10774 ( .A(N5980), .B(n3687), .Z(n2730) );
  CANR2X1 U10775 ( .A(mem_data1[822]), .B(n3898), .C(N9102), .D(n3661), .Z(
        n2729) );
  CND3XL U10776 ( .A(n2732), .B(n2733), .C(n2734), .Z(N10145) );
  CANR2X1 U10777 ( .A(N2897), .B(n3576), .C(n3613), .D(N7458), .Z(n2734) );
  CND2X1 U10778 ( .A(N5979), .B(n3694), .Z(n2733) );
  CANR2X1 U10779 ( .A(mem_data1[821]), .B(n3898), .C(N9101), .D(n3661), .Z(
        n2732) );
  CND3XL U10780 ( .A(n2735), .B(n2736), .C(n2737), .Z(N10144) );
  CANR2X1 U10781 ( .A(N2896), .B(n3576), .C(n3612), .D(N7459), .Z(n2737) );
  CND2X1 U10782 ( .A(N5978), .B(n3697), .Z(n2736) );
  CANR2X1 U10783 ( .A(mem_data1[820]), .B(n3898), .C(N9100), .D(n3661), .Z(
        n2735) );
  CND3XL U10784 ( .A(n2738), .B(n2739), .C(n2740), .Z(N10143) );
  CANR2X1 U10785 ( .A(N2895), .B(n3576), .C(n3612), .D(N7460), .Z(n2740) );
  CND2X1 U10786 ( .A(N5977), .B(n3693), .Z(n2739) );
  CANR2X1 U10787 ( .A(mem_data1[819]), .B(n3898), .C(N9099), .D(n3661), .Z(
        n2738) );
  CND3XL U10788 ( .A(n2741), .B(n2742), .C(n2743), .Z(N10142) );
  CANR2X1 U10789 ( .A(N2894), .B(n3576), .C(n3612), .D(N7461), .Z(n2743) );
  CND2X1 U10790 ( .A(N5976), .B(n3698), .Z(n2742) );
  CANR2X1 U10791 ( .A(mem_data1[818]), .B(n3898), .C(N9098), .D(n3661), .Z(
        n2741) );
  CND3XL U10792 ( .A(n2744), .B(n2745), .C(n2746), .Z(N10141) );
  CANR2X1 U10793 ( .A(N2893), .B(n3576), .C(n3612), .D(N7462), .Z(n2746) );
  CND2X1 U10794 ( .A(N5975), .B(n3689), .Z(n2745) );
  CANR2X1 U10795 ( .A(mem_data1[817]), .B(n3898), .C(N9097), .D(n3661), .Z(
        n2744) );
  CND3XL U10796 ( .A(n2747), .B(n2748), .C(n2749), .Z(N10140) );
  CANR2X1 U10797 ( .A(N2892), .B(n3576), .C(n3612), .D(N7463), .Z(n2749) );
  CND2X1 U10798 ( .A(N5974), .B(n3689), .Z(n2748) );
  CANR2X1 U10799 ( .A(mem_data1[816]), .B(n3898), .C(N9096), .D(n3661), .Z(
        n2747) );
  CND3XL U10800 ( .A(n2750), .B(n2751), .C(n2752), .Z(N10139) );
  CANR2X1 U10801 ( .A(N2891), .B(n3576), .C(n3612), .D(N7464), .Z(n2752) );
  CND2X1 U10802 ( .A(N5973), .B(n3687), .Z(n2751) );
  CANR2X1 U10803 ( .A(mem_data1[815]), .B(n3898), .C(N9095), .D(n3661), .Z(
        n2750) );
  CND3XL U10804 ( .A(n2753), .B(n2754), .C(n2755), .Z(N10138) );
  CANR2X1 U10805 ( .A(N2890), .B(n3576), .C(n3612), .D(N7465), .Z(n2755) );
  CND2X1 U10806 ( .A(N5972), .B(n3688), .Z(n2754) );
  CANR2X1 U10807 ( .A(mem_data1[814]), .B(n3898), .C(N9094), .D(n3661), .Z(
        n2753) );
  CND3XL U10808 ( .A(n2756), .B(n2757), .C(n2758), .Z(N10137) );
  CANR2X1 U10809 ( .A(N2889), .B(n3576), .C(n3612), .D(N7466), .Z(n2758) );
  CND2X1 U10810 ( .A(N5971), .B(n3694), .Z(n2757) );
  CANR2X1 U10811 ( .A(mem_data1[813]), .B(n3898), .C(N9093), .D(n3661), .Z(
        n2756) );
  CND3XL U10812 ( .A(n2759), .B(n2760), .C(n2761), .Z(N10136) );
  CANR2X1 U10813 ( .A(N2888), .B(n3576), .C(n3612), .D(N7467), .Z(n2761) );
  CND2X1 U10814 ( .A(N5970), .B(n3697), .Z(n2760) );
  CANR2X1 U10815 ( .A(mem_data1[812]), .B(n3898), .C(N9092), .D(n3661), .Z(
        n2759) );
  CND3XL U10816 ( .A(n2762), .B(n2763), .C(n2764), .Z(N10135) );
  CANR2X1 U10817 ( .A(N2887), .B(n3578), .C(n3612), .D(N7468), .Z(n2764) );
  CND2X1 U10818 ( .A(N5969), .B(n3690), .Z(n2763) );
  CANR2X1 U10819 ( .A(mem_data1[811]), .B(n3898), .C(N9091), .D(n3661), .Z(
        n2762) );
  CND3XL U10820 ( .A(n2765), .B(n2766), .C(n2767), .Z(N10134) );
  CANR2X1 U10821 ( .A(N2886), .B(n3578), .C(n3612), .D(N7469), .Z(n2767) );
  CND2X1 U10822 ( .A(N5968), .B(n3698), .Z(n2766) );
  CANR2X1 U10823 ( .A(mem_data1[810]), .B(n3898), .C(N9090), .D(n3661), .Z(
        n2765) );
  CND3XL U10824 ( .A(n2768), .B(n2769), .C(n2770), .Z(N10133) );
  CANR2X1 U10825 ( .A(N2885), .B(n3578), .C(n3612), .D(N7470), .Z(n2770) );
  CND2X1 U10826 ( .A(N5967), .B(n3689), .Z(n2769) );
  CANR2X1 U10827 ( .A(mem_data1[809]), .B(n3898), .C(N9089), .D(n3661), .Z(
        n2768) );
  CND3XL U10828 ( .A(n2771), .B(n2772), .C(n2773), .Z(N10132) );
  CANR2X1 U10829 ( .A(N2884), .B(n3578), .C(n3612), .D(N7471), .Z(n2773) );
  CND2X1 U10830 ( .A(N5966), .B(n3688), .Z(n2772) );
  CANR2X1 U10831 ( .A(mem_data1[808]), .B(n3898), .C(N9088), .D(n3661), .Z(
        n2771) );
  CND3XL U10832 ( .A(n2774), .B(n2775), .C(n2776), .Z(N10131) );
  CND3XL U10833 ( .A(n2777), .B(n2778), .C(n2779), .Z(N10130) );
  CND3XL U10834 ( .A(n2780), .B(n2781), .C(n2782), .Z(N10129) );
  CANR2X1 U10835 ( .A(N2881), .B(n3591), .C(n3635), .D(N7474), .Z(n2782) );
  CND2X1 U10836 ( .A(N5963), .B(n3685), .Z(n2781) );
  CANR2X1 U10837 ( .A(mem_data1[805]), .B(n3898), .C(N9085), .D(n3659), .Z(
        n2780) );
  CND3XL U10838 ( .A(n2783), .B(n2784), .C(n2785), .Z(N10128) );
  CANR2X1 U10839 ( .A(N2880), .B(n3591), .C(n3636), .D(N7475), .Z(n2785) );
  CND2X1 U10840 ( .A(N5962), .B(n3684), .Z(n2784) );
  CANR2X1 U10841 ( .A(mem_data1[804]), .B(n3898), .C(N9084), .D(n3659), .Z(
        n2783) );
  CND3XL U10842 ( .A(n2786), .B(n2787), .C(n2788), .Z(N10127) );
  CANR2X1 U10843 ( .A(N2879), .B(n3603), .C(n3636), .D(N7476), .Z(n2788) );
  CND2X1 U10844 ( .A(N5961), .B(n3697), .Z(n2787) );
  CANR2X1 U10845 ( .A(mem_data1[803]), .B(n3898), .C(N9083), .D(n3659), .Z(
        n2786) );
  CND3XL U10846 ( .A(n2789), .B(n2790), .C(n2791), .Z(N10126) );
  CANR2X1 U10847 ( .A(N2878), .B(n3602), .C(n3635), .D(N7477), .Z(n2791) );
  CND2X1 U10848 ( .A(N5960), .B(n3687), .Z(n2790) );
  CANR2X1 U10849 ( .A(mem_data1[802]), .B(n3898), .C(N9082), .D(n3660), .Z(
        n2789) );
  CND3XL U10850 ( .A(n2792), .B(n2793), .C(n2794), .Z(N10125) );
  CANR2X1 U10851 ( .A(N2877), .B(n3602), .C(n3635), .D(N7478), .Z(n2794) );
  CND2X1 U10852 ( .A(N5959), .B(n3688), .Z(n2793) );
  CANR2X1 U10853 ( .A(mem_data1[801]), .B(n3898), .C(N9081), .D(n3660), .Z(
        n2792) );
  CND3XL U10854 ( .A(n2795), .B(n2796), .C(n2797), .Z(N10124) );
  CANR2X1 U10855 ( .A(N2876), .B(n3602), .C(n3635), .D(N7479), .Z(n2797) );
  CND2X1 U10856 ( .A(N5958), .B(n3696), .Z(n2796) );
  CANR2X1 U10857 ( .A(mem_data1[800]), .B(n3898), .C(N9080), .D(n3660), .Z(
        n2795) );
  CND3XL U10858 ( .A(n2798), .B(n2799), .C(n2800), .Z(N10123) );
  CANR2X1 U10859 ( .A(N2875), .B(n3602), .C(n3635), .D(N7480), .Z(n2800) );
  CND2X1 U10860 ( .A(N5957), .B(n3686), .Z(n2799) );
  CANR2X1 U10861 ( .A(mem_data1[799]), .B(n3898), .C(N9079), .D(n3660), .Z(
        n2798) );
  CND3XL U10862 ( .A(n2801), .B(n2802), .C(n2803), .Z(N10122) );
  CANR2X1 U10863 ( .A(N2874), .B(n3602), .C(n3635), .D(N7481), .Z(n2803) );
  CND2X1 U10864 ( .A(N5956), .B(n3698), .Z(n2802) );
  CANR2X1 U10865 ( .A(mem_data1[798]), .B(n3898), .C(N9078), .D(n3660), .Z(
        n2801) );
  CND3XL U10866 ( .A(n2804), .B(n2805), .C(n2806), .Z(N10121) );
  CANR2X1 U10867 ( .A(N2873), .B(n3602), .C(n3635), .D(N7482), .Z(n2806) );
  CND2X1 U10868 ( .A(N5955), .B(n3692), .Z(n2805) );
  CANR2X1 U10869 ( .A(mem_data1[797]), .B(n3898), .C(N9077), .D(n3660), .Z(
        n2804) );
  CND3XL U10870 ( .A(n2807), .B(n2808), .C(n2809), .Z(N10120) );
  CANR2X1 U10871 ( .A(N2872), .B(n3602), .C(n3635), .D(N7483), .Z(n2809) );
  CND2X1 U10872 ( .A(N5954), .B(n3695), .Z(n2808) );
  CANR2X1 U10873 ( .A(mem_data1[796]), .B(n3898), .C(N9076), .D(n3660), .Z(
        n2807) );
  CND3XL U10874 ( .A(n2810), .B(n2811), .C(n2812), .Z(N10119) );
  CANR2X1 U10875 ( .A(N2871), .B(n3602), .C(n3635), .D(N7484), .Z(n2812) );
  CND2X1 U10876 ( .A(N5953), .B(n3692), .Z(n2811) );
  CANR2X1 U10877 ( .A(mem_data1[795]), .B(n3898), .C(N9075), .D(n3660), .Z(
        n2810) );
  CND3XL U10878 ( .A(n2813), .B(n2814), .C(n2815), .Z(N10118) );
  CANR2X1 U10879 ( .A(N2870), .B(n3602), .C(n3626), .D(N7485), .Z(n2815) );
  CND2X1 U10880 ( .A(N5952), .B(n3690), .Z(n2814) );
  CANR2X1 U10881 ( .A(mem_data1[794]), .B(n3898), .C(N9074), .D(n3660), .Z(
        n2813) );
  CND3XL U10882 ( .A(n2816), .B(n2817), .C(n2818), .Z(N10117) );
  CANR2X1 U10883 ( .A(N2869), .B(n3602), .C(n3626), .D(N7486), .Z(n2818) );
  CND2X1 U10884 ( .A(N5951), .B(n3693), .Z(n2817) );
  CANR2X1 U10885 ( .A(mem_data1[793]), .B(n3898), .C(N9073), .D(n3660), .Z(
        n2816) );
  CND3XL U10886 ( .A(n2819), .B(n2820), .C(n2821), .Z(N10116) );
  CANR2X1 U10887 ( .A(N2868), .B(n3602), .C(n3626), .D(N7487), .Z(n2821) );
  CND2X1 U10888 ( .A(N5950), .B(n3683), .Z(n2820) );
  CANR2X1 U10889 ( .A(mem_data1[792]), .B(n3898), .C(N9072), .D(n3660), .Z(
        n2819) );
  CND3XL U10890 ( .A(n2822), .B(n2823), .C(n2824), .Z(N10115) );
  CANR2X1 U10891 ( .A(N2867), .B(n3602), .C(n3626), .D(N7488), .Z(n2824) );
  CND2X1 U10892 ( .A(N5949), .B(n3691), .Z(n2823) );
  CANR2X1 U10893 ( .A(mem_data1[791]), .B(n3898), .C(N9071), .D(n3660), .Z(
        n2822) );
  CND3XL U10894 ( .A(n2825), .B(n2826), .C(n2827), .Z(N10114) );
  CANR2X1 U10895 ( .A(N2866), .B(n3602), .C(n3626), .D(N7489), .Z(n2827) );
  CND2X1 U10896 ( .A(N5948), .B(n3694), .Z(n2826) );
  CANR2X1 U10897 ( .A(mem_data1[790]), .B(n3898), .C(N9070), .D(n3660), .Z(
        n2825) );
  CND3XL U10898 ( .A(n2828), .B(n2829), .C(n2830), .Z(N10113) );
  CANR2X1 U10899 ( .A(N2865), .B(n3602), .C(n3626), .D(N7490), .Z(n2830) );
  CND2X1 U10900 ( .A(N5947), .B(n3689), .Z(n2829) );
  CANR2X1 U10901 ( .A(mem_data1[789]), .B(n3898), .C(N9069), .D(n3660), .Z(
        n2828) );
  CND3XL U10902 ( .A(n2831), .B(n2832), .C(n2833), .Z(N10112) );
  CANR2X1 U10903 ( .A(N2864), .B(n3602), .C(n3626), .D(N7491), .Z(n2833) );
  CND2X1 U10904 ( .A(N5946), .B(n3685), .Z(n2832) );
  CANR2X1 U10905 ( .A(mem_data1[788]), .B(n3898), .C(N9068), .D(n3660), .Z(
        n2831) );
  CND3XL U10906 ( .A(n2834), .B(n2835), .C(n2836), .Z(N10111) );
  CANR2X1 U10907 ( .A(N2863), .B(n3602), .C(n3626), .D(N7492), .Z(n2836) );
  CND2X1 U10908 ( .A(N5945), .B(n3684), .Z(n2835) );
  CANR2X1 U10909 ( .A(mem_data1[787]), .B(n3898), .C(N9067), .D(n3660), .Z(
        n2834) );
  CND3XL U10910 ( .A(n2837), .B(n2838), .C(n2839), .Z(N10110) );
  CANR2X1 U10911 ( .A(N2862), .B(n3602), .C(n3626), .D(N7493), .Z(n2839) );
  CND2X1 U10912 ( .A(N5944), .B(n3697), .Z(n2838) );
  CANR2X1 U10913 ( .A(mem_data1[786]), .B(n3898), .C(N9066), .D(n3660), .Z(
        n2837) );
  CND3XL U10914 ( .A(n2840), .B(n2841), .C(n2842), .Z(N10109) );
  CANR2X1 U10915 ( .A(N2861), .B(n3602), .C(n3626), .D(N7494), .Z(n2842) );
  CND2X1 U10916 ( .A(N5943), .B(n3693), .Z(n2841) );
  CANR2X1 U10917 ( .A(mem_data1[785]), .B(n3898), .C(N9065), .D(n3660), .Z(
        n2840) );
  CND3XL U10918 ( .A(n2843), .B(n2844), .C(n2845), .Z(N10108) );
  CANR2X1 U10919 ( .A(N2860), .B(n3603), .C(n3635), .D(N7495), .Z(n2845) );
  CND2X1 U10920 ( .A(N5942), .B(n3697), .Z(n2844) );
  CANR2X1 U10921 ( .A(mem_data1[784]), .B(n3898), .C(N9064), .D(n3660), .Z(
        n2843) );
  CND3XL U10922 ( .A(n2846), .B(n2847), .C(n2848), .Z(N10107) );
  CANR2X1 U10923 ( .A(N2859), .B(n3603), .C(n3636), .D(N7496), .Z(n2848) );
  CND2X1 U10924 ( .A(N5941), .B(n3683), .Z(n2847) );
  CANR2X1 U10925 ( .A(mem_data1[783]), .B(n3898), .C(N9063), .D(n3669), .Z(
        n2846) );
  CND3XL U10926 ( .A(n2849), .B(n2850), .C(n2851), .Z(N10106) );
  CANR2X1 U10927 ( .A(N2858), .B(n3603), .C(n3636), .D(N7497), .Z(n2851) );
  CND2X1 U10928 ( .A(N5940), .B(n3683), .Z(n2850) );
  CANR2X1 U10929 ( .A(mem_data1[782]), .B(n3898), .C(N9062), .D(n3669), .Z(
        n2849) );
  CND3XL U10930 ( .A(n2852), .B(n2853), .C(n2854), .Z(N10105) );
  CANR2X1 U10931 ( .A(N2857), .B(n3603), .C(n3635), .D(N7498), .Z(n2854) );
  CND2X1 U10932 ( .A(N5939), .B(n3683), .Z(n2853) );
  CANR2X1 U10933 ( .A(mem_data1[781]), .B(n3898), .C(N9061), .D(n3669), .Z(
        n2852) );
  CND3XL U10934 ( .A(n2855), .B(n2856), .C(n2857), .Z(N10104) );
  CANR2X1 U10935 ( .A(N2856), .B(n3602), .C(n3636), .D(N7499), .Z(n2857) );
  CND2X1 U10936 ( .A(N5938), .B(n3683), .Z(n2856) );
  CANR2X1 U10937 ( .A(mem_data1[780]), .B(n3898), .C(N9060), .D(n3669), .Z(
        n2855) );
  CND3XL U10938 ( .A(n2858), .B(n2859), .C(n2860), .Z(N10103) );
  CANR2X1 U10939 ( .A(N2855), .B(n3602), .C(n3636), .D(N7500), .Z(n2860) );
  CND2X1 U10940 ( .A(N5937), .B(n3683), .Z(n2859) );
  CANR2X1 U10941 ( .A(mem_data1[779]), .B(n3898), .C(N9059), .D(n3669), .Z(
        n2858) );
  CND3XL U10942 ( .A(n2861), .B(n2862), .C(n2863), .Z(N10102) );
  CANR2X1 U10943 ( .A(N2854), .B(n3603), .C(n3636), .D(N7501), .Z(n2863) );
  CND2X1 U10944 ( .A(N5936), .B(n3683), .Z(n2862) );
  CANR2X1 U10945 ( .A(mem_data1[778]), .B(n3898), .C(N9058), .D(n3669), .Z(
        n2861) );
  CND3XL U10946 ( .A(n2864), .B(n2865), .C(n2866), .Z(N10101) );
  CANR2X1 U10947 ( .A(N2853), .B(n3603), .C(n3636), .D(N7502), .Z(n2866) );
  CND2X1 U10948 ( .A(N5935), .B(n3683), .Z(n2865) );
  CANR2X1 U10949 ( .A(mem_data1[777]), .B(n3898), .C(N9057), .D(n3669), .Z(
        n2864) );
  CND3XL U10950 ( .A(n2867), .B(n2868), .C(n2869), .Z(N10100) );
  CANR2X1 U10951 ( .A(N2852), .B(n3603), .C(n3636), .D(N7503), .Z(n2869) );
  CND2X1 U10952 ( .A(N5934), .B(n3683), .Z(n2868) );
  CANR2X1 U10953 ( .A(mem_data1[776]), .B(n3898), .C(N9056), .D(n3669), .Z(
        n2867) );
  CND3XL U10954 ( .A(n2870), .B(n2871), .C(n2872), .Z(N10099) );
  CANR2X1 U10955 ( .A(N2851), .B(n3603), .C(n3636), .D(N7504), .Z(n2872) );
  CND2X1 U10956 ( .A(N5933), .B(n3683), .Z(n2871) );
  CANR2X1 U10957 ( .A(mem_data1[775]), .B(n3898), .C(N9055), .D(n3669), .Z(
        n2870) );
  CND3XL U10958 ( .A(n2873), .B(n2874), .C(n2875), .Z(N10098) );
  CANR2X1 U10959 ( .A(N2850), .B(n3603), .C(n3636), .D(N7505), .Z(n2875) );
  CND2X1 U10960 ( .A(N5932), .B(n3683), .Z(n2874) );
  CANR2X1 U10961 ( .A(mem_data1[774]), .B(n3898), .C(N9054), .D(n3669), .Z(
        n2873) );
  CND3XL U10962 ( .A(n2876), .B(n2877), .C(n2878), .Z(N10097) );
  CANR2X1 U10963 ( .A(N2849), .B(n3603), .C(n3637), .D(N7506), .Z(n2878) );
  CND2X1 U10964 ( .A(N5931), .B(n3683), .Z(n2877) );
  CANR2X1 U10965 ( .A(mem_data1[773]), .B(n3898), .C(N9053), .D(n3669), .Z(
        n2876) );
  CND3XL U10966 ( .A(n2879), .B(n2880), .C(n2881), .Z(N10096) );
  CANR2X1 U10967 ( .A(N2848), .B(n3603), .C(n3635), .D(N7507), .Z(n2881) );
  CND2X1 U10968 ( .A(N5930), .B(n3683), .Z(n2880) );
  CANR2X1 U10969 ( .A(mem_data1[772]), .B(n3898), .C(N9052), .D(n3669), .Z(
        n2879) );
  CND3XL U10970 ( .A(n2882), .B(n2883), .C(n2884), .Z(N10095) );
  CANR2X1 U10971 ( .A(N2847), .B(n3603), .C(n3637), .D(N7508), .Z(n2884) );
  CND2X1 U10972 ( .A(N5929), .B(n3683), .Z(n2883) );
  CANR2X1 U10973 ( .A(mem_data1[771]), .B(n3898), .C(N9051), .D(n3669), .Z(
        n2882) );
  CND3XL U10974 ( .A(n2885), .B(n2886), .C(n2887), .Z(N10094) );
  CANR2X1 U10975 ( .A(N2846), .B(n3603), .C(n3636), .D(N7509), .Z(n2887) );
  CND2X1 U10976 ( .A(N5928), .B(n3683), .Z(n2886) );
  CANR2X1 U10977 ( .A(mem_data1[770]), .B(n3898), .C(N9050), .D(n3669), .Z(
        n2885) );
  CND3XL U10978 ( .A(n2888), .B(n2889), .C(n2890), .Z(N10093) );
  CANR2X1 U10979 ( .A(N2845), .B(n3603), .C(n3637), .D(N7510), .Z(n2890) );
  CND2X1 U10980 ( .A(N5927), .B(n3683), .Z(n2889) );
  CANR2X1 U10981 ( .A(mem_data1[769]), .B(n3898), .C(N9049), .D(n3669), .Z(
        n2888) );
  CND3XL U10982 ( .A(n2891), .B(n2892), .C(n2893), .Z(N10092) );
  CANR2X1 U10983 ( .A(N2844), .B(n3603), .C(n3637), .D(N7511), .Z(n2893) );
  CND2X1 U10984 ( .A(N5926), .B(n3683), .Z(n2892) );
  CANR2X1 U10985 ( .A(mem_data1[768]), .B(n3898), .C(N9048), .D(n3669), .Z(
        n2891) );
  CND3XL U10986 ( .A(n2894), .B(n2895), .C(n2896), .Z(N10091) );
  CANR2X1 U10987 ( .A(N2843), .B(n3603), .C(n3637), .D(N7512), .Z(n2896) );
  CND2X1 U10988 ( .A(N5925), .B(n3683), .Z(n2895) );
  CANR2X1 U10989 ( .A(mem_data1[767]), .B(n3898), .C(N9047), .D(n3662), .Z(
        n2894) );
  CND3XL U10990 ( .A(n2897), .B(n2898), .C(n2899), .Z(N10090) );
  CANR2X1 U10991 ( .A(N2842), .B(n3603), .C(n3636), .D(N7513), .Z(n2899) );
  CND2X1 U10992 ( .A(N5924), .B(n3683), .Z(n2898) );
  CANR2X1 U10993 ( .A(mem_data1[766]), .B(n3898), .C(N9046), .D(n3659), .Z(
        n2897) );
  CND3XL U10994 ( .A(n2900), .B(n2901), .C(n2902), .Z(N10089) );
  CANR2X1 U10995 ( .A(N2841), .B(n3603), .C(n3637), .D(N7514), .Z(n2902) );
  CND2X1 U10996 ( .A(N5923), .B(n3683), .Z(n2901) );
  CANR2X1 U10997 ( .A(mem_data1[765]), .B(n3898), .C(N9045), .D(n3659), .Z(
        n2900) );
  CND3XL U10998 ( .A(n2903), .B(n2904), .C(n2905), .Z(N10088) );
  CANR2X1 U10999 ( .A(N2840), .B(n3604), .C(n3636), .D(N7515), .Z(n2905) );
  CND2X1 U11000 ( .A(N5922), .B(n3683), .Z(n2904) );
  CANR2X1 U11001 ( .A(mem_data1[764]), .B(n3898), .C(N9044), .D(n3659), .Z(
        n2903) );
  CND3XL U11002 ( .A(n2906), .B(n2907), .C(n2908), .Z(N10087) );
  CANR2X1 U11003 ( .A(N2839), .B(n3604), .C(n3636), .D(N7516), .Z(n2908) );
  CND2X1 U11004 ( .A(N5921), .B(n3683), .Z(n2907) );
  CANR2X1 U11005 ( .A(mem_data1[763]), .B(n3898), .C(N9043), .D(n3659), .Z(
        n2906) );
  CND3XL U11006 ( .A(n2909), .B(n2910), .C(n2911), .Z(N10086) );
  CANR2X1 U11007 ( .A(N2838), .B(n3603), .C(n3636), .D(N7517), .Z(n2911) );
  CND2X1 U11008 ( .A(N5920), .B(n3687), .Z(n2910) );
  CANR2X1 U11009 ( .A(mem_data1[762]), .B(n3898), .C(N9042), .D(n3659), .Z(
        n2909) );
  CND3XL U11010 ( .A(n2912), .B(n2913), .C(n2914), .Z(N10085) );
  CANR2X1 U11011 ( .A(N2837), .B(n3603), .C(n3636), .D(N7518), .Z(n2914) );
  CND2X1 U11012 ( .A(N5919), .B(n3697), .Z(n2913) );
  CANR2X1 U11013 ( .A(mem_data1[761]), .B(n3898), .C(N9041), .D(n3668), .Z(
        n2912) );
  CND3XL U11014 ( .A(n2915), .B(n2916), .C(n2917), .Z(N10084) );
  CANR2X1 U11015 ( .A(N2836), .B(n3602), .C(n3636), .D(N7519), .Z(n2917) );
  CND2X1 U11016 ( .A(N5918), .B(n3685), .Z(n2916) );
  CANR2X1 U11017 ( .A(mem_data1[760]), .B(n3898), .C(N9040), .D(n3668), .Z(
        n2915) );
  CND3XL U11018 ( .A(n2918), .B(n2919), .C(n2920), .Z(N10083) );
  CANR2X1 U11019 ( .A(N2835), .B(n3603), .C(n3636), .D(N7520), .Z(n2920) );
  CND2X1 U11020 ( .A(N5917), .B(n3698), .Z(n2919) );
  CANR2X1 U11021 ( .A(mem_data1[759]), .B(n3898), .C(N9039), .D(n3668), .Z(
        n2918) );
  CND3XL U11022 ( .A(n2921), .B(n2922), .C(n2923), .Z(N10082) );
  CANR2X1 U11023 ( .A(N2834), .B(n3603), .C(n3636), .D(N7521), .Z(n2923) );
  CND2X1 U11024 ( .A(N5916), .B(n3696), .Z(n2922) );
  CANR2X1 U11025 ( .A(mem_data1[758]), .B(n3898), .C(N9038), .D(n3668), .Z(
        n2921) );
  CND3XL U11026 ( .A(n2924), .B(n2925), .C(n2926), .Z(N10081) );
  CANR2X1 U11027 ( .A(N2833), .B(n3603), .C(n3631), .D(N7522), .Z(n2926) );
  CND2X1 U11028 ( .A(N5915), .B(n3687), .Z(n2925) );
  CANR2X1 U11029 ( .A(mem_data1[757]), .B(n3898), .C(N9037), .D(n3668), .Z(
        n2924) );
  CND3XL U11030 ( .A(n2927), .B(n2928), .C(n2929), .Z(N10080) );
  CANR2X1 U11031 ( .A(N2832), .B(n3602), .C(n3631), .D(N7523), .Z(n2929) );
  CND2X1 U11032 ( .A(N5914), .B(n3698), .Z(n2928) );
  CANR2X1 U11033 ( .A(mem_data1[756]), .B(n3898), .C(N9036), .D(n3668), .Z(
        n2927) );
  CND3XL U11034 ( .A(n2930), .B(n2931), .C(n2932), .Z(N10079) );
  CANR2X1 U11035 ( .A(N2831), .B(n3603), .C(n3631), .D(N7524), .Z(n2932) );
  CND2X1 U11036 ( .A(N5913), .B(n3697), .Z(n2931) );
  CANR2X1 U11037 ( .A(mem_data1[755]), .B(n3898), .C(N9035), .D(n3668), .Z(
        n2930) );
  CND3XL U11038 ( .A(n2933), .B(n2934), .C(n2935), .Z(N10078) );
  CANR2X1 U11039 ( .A(N2830), .B(n3602), .C(n3631), .D(N7525), .Z(n2935) );
  CND2X1 U11040 ( .A(N5912), .B(n3690), .Z(n2934) );
  CANR2X1 U11041 ( .A(mem_data1[754]), .B(n3898), .C(N9034), .D(n3668), .Z(
        n2933) );
  CND3XL U11042 ( .A(n2936), .B(n2937), .C(n2938), .Z(N10077) );
  CANR2X1 U11043 ( .A(N2829), .B(n3597), .C(n3631), .D(N7526), .Z(n2938) );
  CND2X1 U11044 ( .A(N5911), .B(n3697), .Z(n2937) );
  CANR2X1 U11045 ( .A(mem_data1[753]), .B(n3898), .C(N9033), .D(n3668), .Z(
        n2936) );
  CND3XL U11046 ( .A(n2939), .B(n2940), .C(n2941), .Z(N10076) );
  CANR2X1 U11047 ( .A(N2828), .B(n3597), .C(n3631), .D(N7527), .Z(n2941) );
  CND2X1 U11048 ( .A(N5910), .B(n3684), .Z(n2940) );
  CANR2X1 U11049 ( .A(mem_data1[752]), .B(n3898), .C(N9032), .D(n3668), .Z(
        n2939) );
  CND3XL U11050 ( .A(n2942), .B(n2943), .C(n2944), .Z(N10075) );
  CANR2X1 U11051 ( .A(N2827), .B(n3597), .C(n3631), .D(N7528), .Z(n2944) );
  CND2X1 U11052 ( .A(N5909), .B(n3686), .Z(n2943) );
  CANR2X1 U11053 ( .A(mem_data1[751]), .B(n3898), .C(N9031), .D(n3668), .Z(
        n2942) );
  CND3XL U11054 ( .A(n2945), .B(n2946), .C(n2947), .Z(N10074) );
  CANR2X1 U11055 ( .A(N2826), .B(n3597), .C(n3631), .D(N7529), .Z(n2947) );
  CND2X1 U11056 ( .A(N5908), .B(n3688), .Z(n2946) );
  CANR2X1 U11057 ( .A(mem_data1[750]), .B(n3898), .C(N9030), .D(n3668), .Z(
        n2945) );
  CND3XL U11058 ( .A(n2948), .B(n2949), .C(n2950), .Z(N10073) );
  CANR2X1 U11059 ( .A(N2825), .B(n3597), .C(n3631), .D(N7530), .Z(n2950) );
  CND2X1 U11060 ( .A(N5907), .B(n3695), .Z(n2949) );
  CANR2X1 U11061 ( .A(mem_data1[749]), .B(n3898), .C(N9029), .D(n3668), .Z(
        n2948) );
  CND3XL U11062 ( .A(n2951), .B(n2952), .C(n2953), .Z(N10072) );
  CANR2X1 U11063 ( .A(N2824), .B(n3597), .C(n3631), .D(N7531), .Z(n2953) );
  CND2X1 U11064 ( .A(N5906), .B(n3687), .Z(n2952) );
  CANR2X1 U11065 ( .A(mem_data1[748]), .B(n3898), .C(N9028), .D(n3668), .Z(
        n2951) );
  CND3XL U11066 ( .A(n2954), .B(n2955), .C(n2956), .Z(N10071) );
  CANR2X1 U11067 ( .A(N2823), .B(n3597), .C(n3631), .D(N7532), .Z(n2956) );
  CND2X1 U11068 ( .A(N5905), .B(n3686), .Z(n2955) );
  CANR2X1 U11069 ( .A(mem_data1[747]), .B(n3898), .C(N9027), .D(n3668), .Z(
        n2954) );
  CND3XL U11070 ( .A(n2957), .B(n2958), .C(n2959), .Z(N10070) );
  CANR2X1 U11071 ( .A(N2822), .B(n3597), .C(n3631), .D(N7533), .Z(n2959) );
  CND2X1 U11072 ( .A(N5904), .B(n3693), .Z(n2958) );
  CANR2X1 U11073 ( .A(mem_data1[746]), .B(n3898), .C(N9026), .D(n3668), .Z(
        n2957) );
  CND3XL U11074 ( .A(n2960), .B(n2961), .C(n2962), .Z(N10069) );
  CANR2X1 U11075 ( .A(N2821), .B(n3597), .C(n3631), .D(N7534), .Z(n2962) );
  CND2X1 U11076 ( .A(N5903), .B(n3697), .Z(n2961) );
  CANR2X1 U11077 ( .A(mem_data1[745]), .B(n3898), .C(N9025), .D(n3669), .Z(
        n2960) );
  CND3XL U11078 ( .A(n2963), .B(n2964), .C(n2965), .Z(N10068) );
  CANR2X1 U11079 ( .A(N2820), .B(n3597), .C(n3630), .D(N7535), .Z(n2965) );
  CND2X1 U11080 ( .A(N5902), .B(n3688), .Z(n2964) );
  CANR2X1 U11081 ( .A(mem_data1[744]), .B(n3898), .C(N9024), .D(n3669), .Z(
        n2963) );
  CND3XL U11082 ( .A(n2966), .B(n2967), .C(n2968), .Z(N10067) );
  CANR2X1 U11083 ( .A(N2819), .B(n3597), .C(n3630), .D(N7536), .Z(n2968) );
  CND2X1 U11084 ( .A(N5901), .B(n3698), .Z(n2967) );
  CANR2X1 U11085 ( .A(mem_data1[743]), .B(n3898), .C(N9023), .D(n3669), .Z(
        n2966) );
  CND3XL U11086 ( .A(n2969), .B(n2970), .C(n2971), .Z(N10066) );
  CANR2X1 U11087 ( .A(N2818), .B(n3597), .C(n3630), .D(N7537), .Z(n2971) );
  CND2X1 U11088 ( .A(N5900), .B(n3690), .Z(n2970) );
  CANR2X1 U11089 ( .A(mem_data1[742]), .B(n3898), .C(N9022), .D(n3669), .Z(
        n2969) );
  CND3XL U11090 ( .A(n2972), .B(n2973), .C(n2974), .Z(N10065) );
  CANR2X1 U11091 ( .A(N2817), .B(n3597), .C(n3630), .D(N7538), .Z(n2974) );
  CND2X1 U11092 ( .A(N5899), .B(n3690), .Z(n2973) );
  CANR2X1 U11093 ( .A(mem_data1[741]), .B(n3898), .C(N9021), .D(n3669), .Z(
        n2972) );
  CND3XL U11094 ( .A(n2975), .B(n2976), .C(n2977), .Z(N10064) );
  CANR2X1 U11095 ( .A(N2816), .B(n3597), .C(n3630), .D(N7539), .Z(n2977) );
  CND2X1 U11096 ( .A(N5898), .B(n3683), .Z(n2976) );
  CANR2X1 U11097 ( .A(mem_data1[740]), .B(n3898), .C(N9020), .D(n3669), .Z(
        n2975) );
  CND3XL U11098 ( .A(n2978), .B(n2979), .C(n2980), .Z(N10063) );
  CANR2X1 U11099 ( .A(N2815), .B(n3597), .C(n3630), .D(N7540), .Z(n2980) );
  CND2X1 U11100 ( .A(N5897), .B(n3688), .Z(n2979) );
  CANR2X1 U11101 ( .A(mem_data1[739]), .B(n3898), .C(N9019), .D(n3667), .Z(
        n2978) );
  CND3XL U11102 ( .A(n2981), .B(n2982), .C(n2983), .Z(N10062) );
  CANR2X1 U11103 ( .A(N2814), .B(n3597), .C(n3633), .D(N7541), .Z(n2983) );
  CND2X1 U11104 ( .A(N5896), .B(n3694), .Z(n2982) );
  CANR2X1 U11105 ( .A(mem_data1[738]), .B(n3898), .C(N9018), .D(n3667), .Z(
        n2981) );
  CND3XL U11106 ( .A(n2984), .B(n2985), .C(n2986), .Z(N10061) );
  CANR2X1 U11107 ( .A(N2813), .B(n3597), .C(n3635), .D(N7542), .Z(n2986) );
  CND2X1 U11108 ( .A(N5895), .B(n3689), .Z(n2985) );
  CANR2X1 U11109 ( .A(mem_data1[737]), .B(n3898), .C(N9017), .D(n3667), .Z(
        n2984) );
  CND3XL U11110 ( .A(n2987), .B(n2988), .C(n2989), .Z(N10060) );
  CANR2X1 U11111 ( .A(N2812), .B(n3597), .C(n3635), .D(N7543), .Z(n2989) );
  CND2X1 U11112 ( .A(N5894), .B(n3691), .Z(n2988) );
  CANR2X1 U11113 ( .A(mem_data1[736]), .B(n3898), .C(N9016), .D(n3667), .Z(
        n2987) );
  CND3XL U11114 ( .A(n2990), .B(n2991), .C(n2992), .Z(N10059) );
  CANR2X1 U11115 ( .A(N2811), .B(n3597), .C(n3636), .D(N7544), .Z(n2992) );
  CND2X1 U11116 ( .A(N5893), .B(n3695), .Z(n2991) );
  CANR2X1 U11117 ( .A(mem_data1[735]), .B(n3898), .C(N9015), .D(n3667), .Z(
        n2990) );
  CND3XL U11118 ( .A(n2993), .B(n2994), .C(n2995), .Z(N10058) );
  CANR2X1 U11119 ( .A(N2810), .B(n3597), .C(n3636), .D(N7545), .Z(n2995) );
  CND2X1 U11120 ( .A(N5892), .B(n3694), .Z(n2994) );
  CANR2X1 U11121 ( .A(mem_data1[734]), .B(n3898), .C(N9014), .D(n3667), .Z(
        n2993) );
  CND3XL U11122 ( .A(n2996), .B(n2997), .C(n2998), .Z(N10057) );
  CANR2X1 U11123 ( .A(N2809), .B(n3597), .C(n3636), .D(N7546), .Z(n2998) );
  CND2X1 U11124 ( .A(N5891), .B(n3690), .Z(n2997) );
  CANR2X1 U11125 ( .A(mem_data1[733]), .B(n3898), .C(N9013), .D(n3667), .Z(
        n2996) );
  CND3XL U11126 ( .A(n2999), .B(n3000), .C(n3001), .Z(N10056) );
  CANR2X1 U11127 ( .A(N2808), .B(n3596), .C(n3636), .D(N7547), .Z(n3001) );
  CND2X1 U11128 ( .A(N5890), .B(n3695), .Z(n3000) );
  CANR2X1 U11129 ( .A(mem_data1[732]), .B(n3898), .C(N9012), .D(n3667), .Z(
        n2999) );
  CND3XL U11130 ( .A(n3002), .B(n3003), .C(n3004), .Z(N10055) );
  CANR2X1 U11131 ( .A(N2807), .B(n3596), .C(n3632), .D(N7548), .Z(n3004) );
  CND2X1 U11132 ( .A(N5889), .B(n3696), .Z(n3003) );
  CANR2X1 U11133 ( .A(mem_data1[731]), .B(n3898), .C(N9011), .D(n3667), .Z(
        n3002) );
  CND3XL U11134 ( .A(n3005), .B(n3006), .C(n3007), .Z(N10054) );
  CANR2X1 U11135 ( .A(N2806), .B(n3599), .C(n3632), .D(N7549), .Z(n3007) );
  CND2X1 U11136 ( .A(N5888), .B(n3695), .Z(n3006) );
  CANR2X1 U11137 ( .A(mem_data1[730]), .B(n3898), .C(N9010), .D(n3667), .Z(
        n3005) );
  CND3XL U11138 ( .A(n3008), .B(n3009), .C(n3010), .Z(N10053) );
  CANR2X1 U11139 ( .A(N2805), .B(n3598), .C(n3632), .D(N7550), .Z(n3010) );
  CND2X1 U11140 ( .A(N5887), .B(n3690), .Z(n3009) );
  CANR2X1 U11141 ( .A(mem_data1[729]), .B(n3898), .C(N9009), .D(n3667), .Z(
        n3008) );
  CND3XL U11142 ( .A(n3011), .B(n3012), .C(n3013), .Z(N10052) );
  CANR2X1 U11143 ( .A(N2804), .B(n3598), .C(n3632), .D(N7551), .Z(n3013) );
  CND2X1 U11144 ( .A(N5886), .B(n3694), .Z(n3012) );
  CANR2X1 U11145 ( .A(mem_data1[728]), .B(n3898), .C(N9008), .D(n3667), .Z(
        n3011) );
  CND3XL U11146 ( .A(n3014), .B(n3015), .C(n3016), .Z(N10051) );
  CANR2X1 U11147 ( .A(N2803), .B(n3598), .C(n3632), .D(N7552), .Z(n3016) );
  CND2X1 U11148 ( .A(N5885), .B(n3689), .Z(n3015) );
  CANR2X1 U11149 ( .A(mem_data1[727]), .B(n3898), .C(N9007), .D(n3667), .Z(
        n3014) );
  CND3XL U11150 ( .A(n3017), .B(n3018), .C(n3019), .Z(N10050) );
  CANR2X1 U11151 ( .A(N2802), .B(n3598), .C(n3632), .D(N7553), .Z(n3019) );
  CND2X1 U11152 ( .A(N5884), .B(n3691), .Z(n3018) );
  CANR2X1 U11153 ( .A(mem_data1[726]), .B(n3898), .C(N9006), .D(n3667), .Z(
        n3017) );
  CND3XL U11154 ( .A(n3020), .B(n3021), .C(n3022), .Z(N10049) );
  CANR2X1 U11155 ( .A(N2801), .B(n3598), .C(n3632), .D(N7554), .Z(n3022) );
  CND2X1 U11156 ( .A(N5883), .B(n3696), .Z(n3021) );
  CANR2X1 U11157 ( .A(mem_data1[725]), .B(n3898), .C(N9005), .D(n3667), .Z(
        n3020) );
  CND3XL U11158 ( .A(n3023), .B(n3024), .C(n3025), .Z(N10048) );
  CANR2X1 U11159 ( .A(N2800), .B(n3598), .C(n3632), .D(N7555), .Z(n3025) );
  CND2X1 U11160 ( .A(N5882), .B(n3684), .Z(n3024) );
  CANR2X1 U11161 ( .A(mem_data1[724]), .B(n3898), .C(N9004), .D(n3667), .Z(
        n3023) );
  CND3XL U11162 ( .A(n3026), .B(n3027), .C(n3028), .Z(N10047) );
  CANR2X1 U11163 ( .A(N2799), .B(n3598), .C(n3632), .D(N7556), .Z(n3028) );
  CND2X1 U11164 ( .A(N5881), .B(n3696), .Z(n3027) );
  CANR2X1 U11165 ( .A(mem_data1[723]), .B(n3898), .C(N9003), .D(n3668), .Z(
        n3026) );
  CND3XL U11166 ( .A(n3029), .B(n3030), .C(n3031), .Z(N10046) );
  CANR2X1 U11167 ( .A(N2798), .B(n3598), .C(n3632), .D(N7557), .Z(n3031) );
  CND2X1 U11168 ( .A(N5880), .B(n3683), .Z(n3030) );
  CANR2X1 U11169 ( .A(mem_data1[722]), .B(n3898), .C(N9002), .D(n3668), .Z(
        n3029) );
  CND3XL U11170 ( .A(n3032), .B(n3033), .C(n3034), .Z(N10045) );
  CANR2X1 U11171 ( .A(N2797), .B(n3598), .C(n3632), .D(N7558), .Z(n3034) );
  CND2X1 U11172 ( .A(N5879), .B(n3696), .Z(n3033) );
  CANR2X1 U11173 ( .A(mem_data1[721]), .B(n3898), .C(N9001), .D(n3668), .Z(
        n3032) );
  CND3XL U11174 ( .A(n3035), .B(n3036), .C(n3037), .Z(N10044) );
  CANR2X1 U11175 ( .A(N2796), .B(n3598), .C(n3632), .D(N7559), .Z(n3037) );
  CND2X1 U11176 ( .A(N5878), .B(n3695), .Z(n3036) );
  CANR2X1 U11177 ( .A(mem_data1[720]), .B(n3898), .C(N9000), .D(n3668), .Z(
        n3035) );
  CND3XL U11178 ( .A(n3038), .B(n3039), .C(n3040), .Z(N10043) );
  CANR2X1 U11179 ( .A(N2795), .B(n3598), .C(n3632), .D(N7560), .Z(n3040) );
  CND2X1 U11180 ( .A(N5877), .B(n3690), .Z(n3039) );
  CANR2X1 U11181 ( .A(mem_data1[719]), .B(n3898), .C(N8999), .D(n3668), .Z(
        n3038) );
  CND3XL U11182 ( .A(n3041), .B(n3042), .C(n3043), .Z(N10042) );
  CANR2X1 U11183 ( .A(N2794), .B(n3598), .C(n3631), .D(N7561), .Z(n3043) );
  CND2X1 U11184 ( .A(N5876), .B(n3685), .Z(n3042) );
  CANR2X1 U11185 ( .A(mem_data1[718]), .B(n3898), .C(N8998), .D(n3668), .Z(
        n3041) );
  CND3XL U11186 ( .A(n3044), .B(n3045), .C(n3046), .Z(N10041) );
  CANR2X1 U11187 ( .A(N2793), .B(n3598), .C(n3631), .D(N7562), .Z(n3046) );
  CND2X1 U11188 ( .A(N5875), .B(n3687), .Z(n3045) );
  CANR2X1 U11189 ( .A(mem_data1[717]), .B(n3898), .C(N8997), .D(n3666), .Z(
        n3044) );
  CND3XL U11190 ( .A(n3047), .B(n3048), .C(n3049), .Z(N10040) );
  CANR2X1 U11191 ( .A(N2792), .B(n3598), .C(n3631), .D(N7563), .Z(n3049) );
  CND2X1 U11192 ( .A(N5874), .B(n3688), .Z(n3048) );
  CANR2X1 U11193 ( .A(mem_data1[716]), .B(n3898), .C(N8996), .D(n3666), .Z(
        n3047) );
  CND3XL U11194 ( .A(n3050), .B(n3051), .C(n3052), .Z(N10039) );
  CANR2X1 U11195 ( .A(N2791), .B(n3598), .C(n3631), .D(N7564), .Z(n3052) );
  CND2X1 U11196 ( .A(N5873), .B(n3686), .Z(n3051) );
  CANR2X1 U11197 ( .A(mem_data1[715]), .B(n3898), .C(N8995), .D(n3666), .Z(
        n3050) );
  CND3XL U11198 ( .A(n3053), .B(n3054), .C(n3055), .Z(N10038) );
  CANR2X1 U11199 ( .A(N2790), .B(n3598), .C(n3631), .D(N7565), .Z(n3055) );
  CND2X1 U11200 ( .A(N5872), .B(n3698), .Z(n3054) );
  CANR2X1 U11201 ( .A(mem_data1[714]), .B(n3898), .C(N8994), .D(n3666), .Z(
        n3053) );
  CND3XL U11202 ( .A(n3056), .B(n3057), .C(n3058), .Z(N10037) );
  CANR2X1 U11203 ( .A(N2789), .B(n3598), .C(n3631), .D(N7566), .Z(n3058) );
  CND2X1 U11204 ( .A(N5871), .B(n3694), .Z(n3057) );
  CANR2X1 U11205 ( .A(mem_data1[713]), .B(n3898), .C(N8993), .D(n3666), .Z(
        n3056) );
  CND3XL U11206 ( .A(n3059), .B(n3060), .C(n3061), .Z(N10036) );
  CANR2X1 U11207 ( .A(N2788), .B(n3598), .C(n3635), .D(N7567), .Z(n3061) );
  CND2X1 U11208 ( .A(N5870), .B(n3696), .Z(n3060) );
  CANR2X1 U11209 ( .A(mem_data1[712]), .B(n3898), .C(N8992), .D(n3666), .Z(
        n3059) );
  CND3XL U11210 ( .A(n3062), .B(n3063), .C(n3064), .Z(N10035) );
  CANR2X1 U11211 ( .A(N2787), .B(n3598), .C(n3631), .D(N7568), .Z(n3064) );
  CND2X1 U11212 ( .A(N5869), .B(n3688), .Z(n3063) );
  CANR2X1 U11213 ( .A(mem_data1[711]), .B(n3898), .C(N8991), .D(n3666), .Z(
        n3062) );
  CND3XL U11214 ( .A(n3065), .B(n3066), .C(n3067), .Z(N10034) );
  CANR2X1 U11215 ( .A(N2786), .B(n3598), .C(n3631), .D(N7569), .Z(n3067) );
  CND2X1 U11216 ( .A(N5868), .B(n3689), .Z(n3066) );
  CANR2X1 U11217 ( .A(mem_data1[710]), .B(n3898), .C(N8990), .D(n3666), .Z(
        n3065) );
  CND3XL U11218 ( .A(n3068), .B(n3069), .C(n3070), .Z(N10033) );
  CANR2X1 U11219 ( .A(N2785), .B(n3598), .C(n3631), .D(N7570), .Z(n3070) );
  CND2X1 U11220 ( .A(N5867), .B(n3693), .Z(n3069) );
  CANR2X1 U11221 ( .A(mem_data1[709]), .B(n3898), .C(N8989), .D(n3666), .Z(
        n3068) );
  CND3XL U11222 ( .A(n3071), .B(n3072), .C(n3073), .Z(N10032) );
  CANR2X1 U11223 ( .A(N2784), .B(n3598), .C(n3631), .D(N7571), .Z(n3073) );
  CND2X1 U11224 ( .A(N5866), .B(n3683), .Z(n3072) );
  CANR2X1 U11225 ( .A(mem_data1[708]), .B(n3898), .C(N8988), .D(n3666), .Z(
        n3071) );
  CND3XL U11226 ( .A(n3074), .B(n3075), .C(n3076), .Z(N10031) );
  CANR2X1 U11227 ( .A(N2783), .B(n3602), .C(n3631), .D(N7572), .Z(n3076) );
  CND2X1 U11228 ( .A(N5865), .B(n3688), .Z(n3075) );
  CANR2X1 U11229 ( .A(mem_data1[707]), .B(n3898), .C(N8987), .D(n3666), .Z(
        n3074) );
  CND3XL U11230 ( .A(n3077), .B(n3078), .C(n3079), .Z(N10030) );
  CANR2X1 U11231 ( .A(N2782), .B(n3597), .C(n3631), .D(N7573), .Z(n3079) );
  CND2X1 U11232 ( .A(N5864), .B(n3691), .Z(n3078) );
  CANR2X1 U11233 ( .A(mem_data1[706]), .B(n3898), .C(N8986), .D(n3666), .Z(
        n3077) );
  CND3XL U11234 ( .A(n3080), .B(n3081), .C(n3082), .Z(N10029) );
  CANR2X1 U11235 ( .A(N2781), .B(n3597), .C(n3631), .D(N7574), .Z(n3082) );
  CND2X1 U11236 ( .A(N5863), .B(n3687), .Z(n3081) );
  CANR2X1 U11237 ( .A(mem_data1[705]), .B(n3898), .C(N8985), .D(n3666), .Z(
        n3080) );
  CND3XL U11238 ( .A(n3083), .B(n3084), .C(n3085), .Z(N10028) );
  CANR2X1 U11239 ( .A(N2780), .B(n3599), .C(n3633), .D(N7575), .Z(n3085) );
  CND2X1 U11240 ( .A(N5862), .B(n3687), .Z(n3084) );
  CANR2X1 U11241 ( .A(mem_data1[704]), .B(n3898), .C(N8984), .D(n3666), .Z(
        n3083) );
  CND3XL U11242 ( .A(n3086), .B(n3087), .C(n3088), .Z(N10027) );
  CANR2X1 U11243 ( .A(N2779), .B(n3599), .C(n3633), .D(N7576), .Z(n3088) );
  CND2X1 U11244 ( .A(N5861), .B(n3687), .Z(n3087) );
  CANR2X1 U11245 ( .A(mem_data1[703]), .B(n3898), .C(N8983), .D(n3666), .Z(
        n3086) );
  CND3XL U11246 ( .A(n3089), .B(n3090), .C(n3091), .Z(N10026) );
  CANR2X1 U11247 ( .A(N2778), .B(n3599), .C(n3633), .D(N7577), .Z(n3091) );
  CND2X1 U11248 ( .A(N5860), .B(n3687), .Z(n3090) );
  CANR2X1 U11249 ( .A(mem_data1[702]), .B(n3898), .C(N8982), .D(n3666), .Z(
        n3089) );
  CND3XL U11250 ( .A(n3092), .B(n3093), .C(n3094), .Z(N10025) );
  CANR2X1 U11251 ( .A(N2777), .B(n3599), .C(n3633), .D(N7578), .Z(n3094) );
  CND2X1 U11252 ( .A(N5859), .B(n3687), .Z(n3093) );
  CANR2X1 U11253 ( .A(mem_data1[701]), .B(n3898), .C(N8981), .D(n3666), .Z(
        n3092) );
  CND3XL U11254 ( .A(n3095), .B(n3096), .C(n3097), .Z(N10024) );
  CANR2X1 U11255 ( .A(N2776), .B(n3599), .C(n3633), .D(N7579), .Z(n3097) );
  CND2X1 U11256 ( .A(N5858), .B(n3687), .Z(n3096) );
  CANR2X1 U11257 ( .A(mem_data1[700]), .B(n3898), .C(N8980), .D(n3667), .Z(
        n3095) );
  CND3XL U11258 ( .A(n3098), .B(n3099), .C(n3100), .Z(N10023) );
  CANR2X1 U11259 ( .A(N2775), .B(n3599), .C(n3633), .D(N7580), .Z(n3100) );
  CND2X1 U11260 ( .A(N5857), .B(n3687), .Z(n3099) );
  CANR2X1 U11261 ( .A(mem_data1[699]), .B(n3898), .C(N8979), .D(n3667), .Z(
        n3098) );
  CND3XL U11262 ( .A(n3101), .B(n3102), .C(n3103), .Z(N10022) );
  CANR2X1 U11263 ( .A(N2774), .B(n3599), .C(n3633), .D(N7581), .Z(n3103) );
  CND2X1 U11264 ( .A(N5856), .B(n3687), .Z(n3102) );
  CANR2X1 U11265 ( .A(mem_data1[698]), .B(n3898), .C(N8978), .D(n3667), .Z(
        n3101) );
  CND3XL U11266 ( .A(n3104), .B(n3105), .C(n3106), .Z(N10021) );
  CANR2X1 U11267 ( .A(N2773), .B(n3599), .C(n3633), .D(N7582), .Z(n3106) );
  CND2X1 U11268 ( .A(N5855), .B(n3687), .Z(n3105) );
  CANR2X1 U11269 ( .A(mem_data1[697]), .B(n3898), .C(N8977), .D(n3667), .Z(
        n3104) );
  CND3XL U11270 ( .A(n3107), .B(n3108), .C(n3109), .Z(N10020) );
  CANR2X1 U11271 ( .A(N2772), .B(n3599), .C(n3633), .D(N7583), .Z(n3109) );
  CND2X1 U11272 ( .A(N5854), .B(n3687), .Z(n3108) );
  CANR2X1 U11273 ( .A(mem_data1[696]), .B(n3898), .C(N8976), .D(n3667), .Z(
        n3107) );
  CND3XL U11274 ( .A(n3110), .B(n3111), .C(n3112), .Z(N10019) );
  CANR2X1 U11275 ( .A(N2771), .B(n3599), .C(n3633), .D(N7584), .Z(n3112) );
  CND2X1 U11276 ( .A(N5853), .B(n3684), .Z(n3111) );
  CANR2X1 U11277 ( .A(mem_data1[695]), .B(n3898), .C(N8975), .D(n3648), .Z(
        n3110) );
  CND3XL U11278 ( .A(n3113), .B(n3114), .C(n3115), .Z(N10018) );
  CANR2X1 U11279 ( .A(N2770), .B(n3599), .C(n3633), .D(N7585), .Z(n3115) );
  CND2X1 U11280 ( .A(N5852), .B(n3691), .Z(n3114) );
  CANR2X1 U11281 ( .A(mem_data1[694]), .B(n3898), .C(N8974), .D(n3670), .Z(
        n3113) );
  CND3XL U11282 ( .A(n3116), .B(n3117), .C(n3118), .Z(N10017) );
  CANR2X1 U11283 ( .A(N2769), .B(n3599), .C(n3633), .D(N7586), .Z(n3118) );
  CND2X1 U11284 ( .A(N5851), .B(n3687), .Z(n3117) );
  CANR2X1 U11285 ( .A(mem_data1[693]), .B(n3898), .C(N8973), .D(n3667), .Z(
        n3116) );
  CND3XL U11286 ( .A(n3119), .B(n3120), .C(n3121), .Z(N10016) );
  CANR2X1 U11287 ( .A(N2768), .B(n3599), .C(n3633), .D(N7587), .Z(n3121) );
  CND2X1 U11288 ( .A(N5850), .B(n3696), .Z(n3120) );
  CANR2X1 U11289 ( .A(mem_data1[692]), .B(n3898), .C(N8972), .D(n3664), .Z(
        n3119) );
  CND3XL U11290 ( .A(n3122), .B(n3123), .C(n3124), .Z(N10015) );
  CANR2X1 U11291 ( .A(N2767), .B(n3599), .C(n3632), .D(N7588), .Z(n3124) );
  CND2X1 U11292 ( .A(N5849), .B(n3698), .Z(n3123) );
  CANR2X1 U11293 ( .A(mem_data1[691]), .B(n3898), .C(N8971), .D(n3664), .Z(
        n3122) );
  CND3XL U11294 ( .A(n3125), .B(n3126), .C(n3127), .Z(N10014) );
  CANR2X1 U11295 ( .A(N2766), .B(n3599), .C(n3632), .D(N7589), .Z(n3127) );
  CND2X1 U11296 ( .A(N5848), .B(n3692), .Z(n3126) );
  CANR2X1 U11297 ( .A(mem_data1[690]), .B(n3898), .C(N8970), .D(n3664), .Z(
        n3125) );
  CND3XL U11298 ( .A(n3128), .B(n3129), .C(n3130), .Z(N10013) );
  CANR2X1 U11299 ( .A(N2765), .B(n3599), .C(n3632), .D(N7590), .Z(n3130) );
  CND2X1 U11300 ( .A(N5847), .B(n3690), .Z(n3129) );
  CANR2X1 U11301 ( .A(mem_data1[689]), .B(n3898), .C(N8969), .D(n3664), .Z(
        n3128) );
  CND3XL U11302 ( .A(n3131), .B(n3132), .C(n3133), .Z(N10012) );
  CANR2X1 U11303 ( .A(N2764), .B(n3599), .C(n3632), .D(N7591), .Z(n3133) );
  CND2X1 U11304 ( .A(N5846), .B(n3686), .Z(n3132) );
  CANR2X1 U11305 ( .A(mem_data1[688]), .B(n3898), .C(N8968), .D(n3665), .Z(
        n3131) );
  CND3XL U11306 ( .A(n3134), .B(n3135), .C(n3136), .Z(N10011) );
  CND3XL U11307 ( .A(n3137), .B(n3138), .C(n3139), .Z(N10010) );
  CND3XL U11308 ( .A(n3140), .B(n3141), .C(n3142), .Z(N10009) );
  CND3XL U11309 ( .A(n3143), .B(n3144), .C(n3145), .Z(N10008) );
  CND3XL U11310 ( .A(n3146), .B(n3147), .C(n3148), .Z(N10007) );
  CND3XL U11311 ( .A(n3149), .B(n3150), .C(n3151), .Z(N10006) );
  CND3XL U11312 ( .A(n3152), .B(n3153), .C(n3154), .Z(N10005) );
  CND3XL U11313 ( .A(n3155), .B(n3156), .C(n3157), .Z(N10004) );
  CND3XL U11314 ( .A(n3158), .B(n3159), .C(n3160), .Z(N10003) );
  CND3XL U11315 ( .A(n3161), .B(n3162), .C(n3163), .Z(N10002) );
  CND3XL U11316 ( .A(n3164), .B(n3165), .C(n3166), .Z(N10001) );
  CND3XL U11317 ( .A(n76), .B(n77), .C(n78), .Z(N9999) );
  CND3XL U11318 ( .A(n80), .B(n81), .C(n82), .Z(N9998) );
  CND3XL U11319 ( .A(n83), .B(n84), .C(n85), .Z(N9997) );
  CND3XL U11320 ( .A(n86), .B(n87), .C(n88), .Z(N9996) );
  CANR2X1 U11321 ( .A(N2748), .B(n3572), .C(n3608), .D(N7607), .Z(n88) );
  CND3XL U11322 ( .A(n89), .B(n90), .C(n91), .Z(N9995) );
  CND3XL U11323 ( .A(n92), .B(n93), .C(n94), .Z(N9994) );
  CND3XL U11324 ( .A(n95), .B(n96), .C(n97), .Z(N9993) );
  CND3XL U11325 ( .A(n98), .B(n99), .C(n100), .Z(N9992) );
  CND3XL U11326 ( .A(n101), .B(n102), .C(n103), .Z(N9991) );
  CND3XL U11327 ( .A(n104), .B(n105), .C(n106), .Z(N9990) );
  CANR2X1 U11328 ( .A(N2742), .B(n3572), .C(n3607), .D(N7613), .Z(n106) );
  CND2X1 U11329 ( .A(N5824), .B(n3687), .Z(n105) );
  CANR2X1 U11330 ( .A(mem_data1[666]), .B(n3898), .C(N8946), .D(n3666), .Z(
        n104) );
  CND3XL U11331 ( .A(n107), .B(n108), .C(n109), .Z(N9989) );
  CANR2X1 U11332 ( .A(N2741), .B(n3572), .C(n3607), .D(N7614), .Z(n109) );
  CND2X1 U11333 ( .A(N5823), .B(n3687), .Z(n108) );
  CANR2X1 U11334 ( .A(mem_data1[665]), .B(n3898), .C(N8945), .D(n3666), .Z(
        n107) );
  CND3XL U11335 ( .A(n110), .B(n111), .C(n112), .Z(N9988) );
  CANR2X1 U11336 ( .A(N2740), .B(n3572), .C(n3607), .D(N7615), .Z(n112) );
  CND2X1 U11337 ( .A(N5822), .B(n3687), .Z(n111) );
  CANR2X1 U11338 ( .A(mem_data1[664]), .B(n3898), .C(N8944), .D(n3666), .Z(
        n110) );
  CND3XL U11339 ( .A(n113), .B(n114), .C(n115), .Z(N9987) );
  CANR2X1 U11340 ( .A(N2739), .B(n3572), .C(n3607), .D(N7616), .Z(n115) );
  CND2X1 U11341 ( .A(N5821), .B(n3689), .Z(n114) );
  CANR2X1 U11342 ( .A(mem_data1[663]), .B(n3898), .C(N8943), .D(n3666), .Z(
        n113) );
  CND3XL U11343 ( .A(n116), .B(n117), .C(n118), .Z(N9986) );
  CANR2X1 U11344 ( .A(N2738), .B(n3572), .C(n3609), .D(N7617), .Z(n118) );
  CND2X1 U11345 ( .A(N5820), .B(n3683), .Z(n117) );
  CANR2X1 U11346 ( .A(mem_data1[662]), .B(n3898), .C(N8942), .D(n3666), .Z(
        n116) );
  CND3XL U11347 ( .A(n119), .B(n120), .C(n121), .Z(N9985) );
  CANR2X1 U11348 ( .A(N2737), .B(n3571), .C(n3609), .D(N7618), .Z(n121) );
  CND2X1 U11349 ( .A(N5819), .B(n3697), .Z(n120) );
  CANR2X1 U11350 ( .A(mem_data1[661]), .B(n3898), .C(N8941), .D(n3652), .Z(
        n119) );
  CND3XL U11351 ( .A(n122), .B(n123), .C(n124), .Z(N9984) );
  CANR2X1 U11352 ( .A(N2736), .B(n3573), .C(n3609), .D(N7619), .Z(n124) );
  CND2X1 U11353 ( .A(N5818), .B(n3687), .Z(n123) );
  CANR2X1 U11354 ( .A(mem_data1[660]), .B(n3898), .C(N8940), .D(n3652), .Z(
        n122) );
  CND3XL U11355 ( .A(n125), .B(n126), .C(n127), .Z(N9983) );
  CANR2X1 U11356 ( .A(N2735), .B(n3573), .C(n3609), .D(N7620), .Z(n127) );
  CND2X1 U11357 ( .A(N5817), .B(n3688), .Z(n126) );
  CANR2X1 U11358 ( .A(mem_data1[659]), .B(n3898), .C(N8939), .D(n3652), .Z(
        n125) );
  CND3XL U11359 ( .A(n128), .B(n129), .C(n130), .Z(N9982) );
  CANR2X1 U11360 ( .A(N2734), .B(n3573), .C(n3609), .D(N7621), .Z(n130) );
  CND2X1 U11361 ( .A(N5816), .B(n3686), .Z(n129) );
  CANR2X1 U11362 ( .A(mem_data1[658]), .B(n3898), .C(N8938), .D(n3652), .Z(
        n128) );
  CND3XL U11363 ( .A(n131), .B(n132), .C(n133), .Z(N9981) );
  CANR2X1 U11364 ( .A(N2733), .B(n3573), .C(n3609), .D(N7622), .Z(n133) );
  CND2X1 U11365 ( .A(N5815), .B(n3698), .Z(n132) );
  CANR2X1 U11366 ( .A(mem_data1[657]), .B(n3898), .C(N8937), .D(n3652), .Z(
        n131) );
  CND3XL U11367 ( .A(n134), .B(n135), .C(n136), .Z(N9980) );
  CANR2X1 U11368 ( .A(N2732), .B(n3573), .C(n3609), .D(N7623), .Z(n136) );
  CND2X1 U11369 ( .A(N5814), .B(n3695), .Z(n135) );
  CANR2X1 U11370 ( .A(mem_data1[656]), .B(n3898), .C(N8936), .D(n3652), .Z(
        n134) );
  CND3XL U11371 ( .A(n137), .B(n138), .C(n139), .Z(N9979) );
  CANR2X1 U11372 ( .A(N2731), .B(n3573), .C(n3609), .D(N7624), .Z(n139) );
  CND2X1 U11373 ( .A(N5813), .B(n3695), .Z(n138) );
  CANR2X1 U11374 ( .A(mem_data1[655]), .B(n3898), .C(N8935), .D(n3652), .Z(
        n137) );
  CND3XL U11375 ( .A(n140), .B(n141), .C(n142), .Z(N9978) );
  CANR2X1 U11376 ( .A(N2730), .B(n3573), .C(n3608), .D(N7625), .Z(n142) );
  CND2X1 U11377 ( .A(N5812), .B(n3693), .Z(n141) );
  CANR2X1 U11378 ( .A(mem_data1[654]), .B(n3898), .C(N8934), .D(n3652), .Z(
        n140) );
  CND3XL U11379 ( .A(n143), .B(n144), .C(n145), .Z(N9977) );
  CANR2X1 U11380 ( .A(N2729), .B(n3573), .C(n3608), .D(N7626), .Z(n145) );
  CND2X1 U11381 ( .A(N5811), .B(n3692), .Z(n144) );
  CANR2X1 U11382 ( .A(mem_data1[653]), .B(n3898), .C(N8933), .D(n3652), .Z(
        n143) );
  CND3XL U11383 ( .A(n146), .B(n147), .C(n148), .Z(N9976) );
  CANR2X1 U11384 ( .A(N2728), .B(n3573), .C(n3608), .D(N7627), .Z(n148) );
  CND2X1 U11385 ( .A(N5810), .B(n3683), .Z(n147) );
  CANR2X1 U11386 ( .A(mem_data1[652]), .B(n3898), .C(N8932), .D(n3652), .Z(
        n146) );
  CND3XL U11387 ( .A(n149), .B(n150), .C(n151), .Z(N9975) );
  CANR2X1 U11388 ( .A(N2727), .B(n3573), .C(n3608), .D(N7628), .Z(n151) );
  CND2X1 U11389 ( .A(N5809), .B(n3694), .Z(n150) );
  CANR2X1 U11390 ( .A(mem_data1[651]), .B(n3898), .C(N8931), .D(n3652), .Z(
        n149) );
  CND3XL U11391 ( .A(n152), .B(n153), .C(n154), .Z(N9974) );
  CANR2X1 U11392 ( .A(N2726), .B(n3573), .C(n3608), .D(N7629), .Z(n154) );
  CND2X1 U11393 ( .A(N5808), .B(n3690), .Z(n153) );
  CANR2X1 U11394 ( .A(mem_data1[650]), .B(n3898), .C(N8930), .D(n3652), .Z(
        n152) );
  CND3XL U11395 ( .A(n155), .B(n156), .C(n157), .Z(N9973) );
  CANR2X1 U11396 ( .A(N2725), .B(n3573), .C(n3608), .D(N7630), .Z(n157) );
  CND2X1 U11397 ( .A(N5807), .B(n3685), .Z(n156) );
  CANR2X1 U11398 ( .A(mem_data1[649]), .B(n3898), .C(N8929), .D(n3652), .Z(
        n155) );
  CND3XL U11399 ( .A(n158), .B(n159), .C(n160), .Z(N9972) );
  CANR2X1 U11400 ( .A(N2724), .B(n3573), .C(n3608), .D(N7631), .Z(n160) );
  CND2X1 U11401 ( .A(N5806), .B(n3696), .Z(n159) );
  CANR2X1 U11402 ( .A(mem_data1[648]), .B(n3898), .C(N8928), .D(n3652), .Z(
        n158) );
  CND3XL U11403 ( .A(n161), .B(n162), .C(n163), .Z(N9971) );
  CANR2X1 U11404 ( .A(N2723), .B(n3573), .C(n3608), .D(N7632), .Z(n163) );
  CND2X1 U11405 ( .A(N5805), .B(n3692), .Z(n162) );
  CANR2X1 U11406 ( .A(mem_data1[647]), .B(n3898), .C(N8927), .D(n3652), .Z(
        n161) );
  CND3XL U11407 ( .A(n164), .B(n165), .C(n166), .Z(N9970) );
  CANR2X1 U11408 ( .A(N2722), .B(n3573), .C(n3608), .D(N7633), .Z(n166) );
  CND2X1 U11409 ( .A(N5804), .B(n3695), .Z(n165) );
  CANR2X1 U11410 ( .A(mem_data1[646]), .B(n3898), .C(N8926), .D(n3651), .Z(
        n164) );
  CND3XL U11411 ( .A(n167), .B(n168), .C(n169), .Z(N9969) );
  CND3XL U11412 ( .A(n170), .B(n171), .C(n172), .Z(N9968) );
  CND3XL U11413 ( .A(n173), .B(n174), .C(n175), .Z(N9967) );
  CND3XL U11414 ( .A(n176), .B(n177), .C(n178), .Z(N9966) );
  CND2X1 U11415 ( .A(N5800), .B(n3684), .Z(n177) );
  CND3XL U11416 ( .A(n179), .B(n180), .C(n181), .Z(N9965) );
  CANR2X1 U11417 ( .A(N2717), .B(n3572), .C(n3608), .D(N7638), .Z(n181) );
  CND2X1 U11418 ( .A(N5799), .B(n3697), .Z(n180) );
  CANR2X1 U11419 ( .A(mem_data1[641]), .B(n3898), .C(N8921), .D(n3655), .Z(
        n179) );
  CND3XL U11420 ( .A(n182), .B(n183), .C(n184), .Z(N9964) );
  CANR2X1 U11421 ( .A(N2716), .B(n3572), .C(n3608), .D(N7639), .Z(n184) );
  CND2X1 U11422 ( .A(N5798), .B(n3686), .Z(n183) );
  CANR2X1 U11423 ( .A(mem_data1[640]), .B(n3898), .C(N8920), .D(n3659), .Z(
        n182) );
  CND3XL U11424 ( .A(n185), .B(n186), .C(n187), .Z(N9963) );
  CANR2X1 U11425 ( .A(N2715), .B(n3572), .C(n3608), .D(N7640), .Z(n187) );
  CND2X1 U11426 ( .A(N5797), .B(n3688), .Z(n186) );
  CANR2X1 U11427 ( .A(mem_data1[639]), .B(n3898), .C(N8919), .D(n3653), .Z(
        n185) );
  CND3XL U11428 ( .A(n188), .B(n189), .C(n190), .Z(N9962) );
  CANR2X1 U11429 ( .A(N2714), .B(n3572), .C(n3608), .D(N7641), .Z(n190) );
  CND2X1 U11430 ( .A(N5796), .B(n3688), .Z(n189) );
  CANR2X1 U11431 ( .A(mem_data1[638]), .B(n3898), .C(N8918), .D(n3653), .Z(
        n188) );
  CND3XL U11432 ( .A(n191), .B(n192), .C(n193), .Z(N9961) );
  CANR2X1 U11433 ( .A(N2713), .B(n3572), .C(n3608), .D(N7642), .Z(n193) );
  CND2X1 U11434 ( .A(N5795), .B(n3688), .Z(n192) );
  CANR2X1 U11435 ( .A(mem_data1[637]), .B(n3898), .C(N8917), .D(n3653), .Z(
        n191) );
  CND3XL U11436 ( .A(n194), .B(n195), .C(n196), .Z(N9960) );
  CANR2X1 U11437 ( .A(N2712), .B(n3572), .C(n3608), .D(N7643), .Z(n196) );
  CND2X1 U11438 ( .A(N5794), .B(n3688), .Z(n195) );
  CANR2X1 U11439 ( .A(mem_data1[636]), .B(n3898), .C(N8916), .D(n3653), .Z(
        n194) );
  CND3XL U11440 ( .A(n197), .B(n198), .C(n199), .Z(N9959) );
  CANR2X1 U11441 ( .A(N2711), .B(n3583), .C(n3618), .D(N7644), .Z(n199) );
  CND2X1 U11442 ( .A(N5793), .B(n3688), .Z(n198) );
  CANR2X1 U11443 ( .A(mem_data1[635]), .B(n3898), .C(N8915), .D(n3653), .Z(
        n197) );
  CND3XL U11444 ( .A(n200), .B(n201), .C(n202), .Z(N9958) );
  CANR2X1 U11445 ( .A(N2710), .B(n3583), .C(n3618), .D(N7645), .Z(n202) );
  CND2X1 U11446 ( .A(N5792), .B(n3688), .Z(n201) );
  CANR2X1 U11447 ( .A(mem_data1[634]), .B(n3898), .C(N8914), .D(n3653), .Z(
        n200) );
  CND3XL U11448 ( .A(n203), .B(n204), .C(n205), .Z(N9957) );
  CANR2X1 U11449 ( .A(N2709), .B(n3585), .C(n3618), .D(N7646), .Z(n205) );
  CND2X1 U11450 ( .A(N5791), .B(n3688), .Z(n204) );
  CANR2X1 U11451 ( .A(mem_data1[633]), .B(n3898), .C(N8913), .D(n3653), .Z(
        n203) );
  CND3XL U11452 ( .A(n206), .B(n207), .C(n208), .Z(N9956) );
  CANR2X1 U11453 ( .A(N2708), .B(n3574), .C(n3620), .D(N7647), .Z(n208) );
  CND2X1 U11454 ( .A(N5790), .B(n3688), .Z(n207) );
  CANR2X1 U11455 ( .A(mem_data1[632]), .B(n3898), .C(N8912), .D(n3653), .Z(
        n206) );
  CND3XL U11456 ( .A(n209), .B(n210), .C(n211), .Z(N9955) );
  CANR2X1 U11457 ( .A(N2707), .B(n3574), .C(n3610), .D(N7648), .Z(n211) );
  CND2X1 U11458 ( .A(N5789), .B(n3688), .Z(n210) );
  CANR2X1 U11459 ( .A(mem_data1[631]), .B(n3898), .C(N8911), .D(n3653), .Z(
        n209) );
  CND3XL U11460 ( .A(n212), .B(n213), .C(n214), .Z(N9954) );
  CANR2X1 U11461 ( .A(N2706), .B(n3574), .C(n3610), .D(N7649), .Z(n214) );
  CND2X1 U11462 ( .A(N5788), .B(n3688), .Z(n213) );
  CANR2X1 U11463 ( .A(mem_data1[630]), .B(n3898), .C(N8910), .D(n3653), .Z(
        n212) );
  CND3XL U11464 ( .A(n215), .B(n216), .C(n217), .Z(N9953) );
  CANR2X1 U11465 ( .A(N2705), .B(n3574), .C(n3610), .D(N7650), .Z(n217) );
  CND2X1 U11466 ( .A(N5787), .B(n3688), .Z(n216) );
  CANR2X1 U11467 ( .A(mem_data1[629]), .B(n3898), .C(N8909), .D(n3653), .Z(
        n215) );
  CND3XL U11468 ( .A(n218), .B(n219), .C(n220), .Z(N9952) );
  CANR2X1 U11469 ( .A(N2704), .B(n3574), .C(n3610), .D(N7651), .Z(n220) );
  CND2X1 U11470 ( .A(N5786), .B(n3696), .Z(n219) );
  CANR2X1 U11471 ( .A(mem_data1[628]), .B(n3898), .C(N8908), .D(n3653), .Z(
        n218) );
  CND3XL U11472 ( .A(n221), .B(n222), .C(n223), .Z(N9951) );
  CANR2X1 U11473 ( .A(N2703), .B(n3574), .C(n3609), .D(N7652), .Z(n223) );
  CND2X1 U11474 ( .A(N5785), .B(n3685), .Z(n222) );
  CANR2X1 U11475 ( .A(mem_data1[627]), .B(n3898), .C(N8907), .D(n3653), .Z(
        n221) );
  CND3XL U11476 ( .A(n224), .B(n225), .C(n226), .Z(N9950) );
  CANR2X1 U11477 ( .A(N2702), .B(n3574), .C(n3609), .D(N7653), .Z(n226) );
  CND2X1 U11478 ( .A(N5784), .B(n3689), .Z(n225) );
  CANR2X1 U11479 ( .A(mem_data1[626]), .B(n3898), .C(N8906), .D(n3653), .Z(
        n224) );
  CND3XL U11480 ( .A(n227), .B(n228), .C(n229), .Z(N9949) );
  CANR2X1 U11481 ( .A(N2701), .B(n3574), .C(n3609), .D(N7654), .Z(n229) );
  CND2X1 U11482 ( .A(N5783), .B(n3691), .Z(n228) );
  CANR2X1 U11483 ( .A(mem_data1[625]), .B(n3898), .C(N8905), .D(n3653), .Z(
        n227) );
  CND3XL U11484 ( .A(n230), .B(n231), .C(n232), .Z(N9948) );
  CANR2X1 U11485 ( .A(N2700), .B(n3574), .C(n3609), .D(N7655), .Z(n232) );
  CND2X1 U11486 ( .A(N5782), .B(n3690), .Z(n231) );
  CANR2X1 U11487 ( .A(mem_data1[624]), .B(n3898), .C(N8904), .D(n3652), .Z(
        n230) );
  CND3XL U11488 ( .A(n233), .B(n234), .C(n235), .Z(N9947) );
  CANR2X1 U11489 ( .A(N2699), .B(n3574), .C(n3609), .D(N7656), .Z(n235) );
  CND2X1 U11490 ( .A(N5781), .B(n3684), .Z(n234) );
  CANR2X1 U11491 ( .A(mem_data1[623]), .B(n3898), .C(N8903), .D(n3652), .Z(
        n233) );
  CND3XL U11492 ( .A(n236), .B(n237), .C(n238), .Z(N9946) );
  CANR2X1 U11493 ( .A(N2698), .B(n3574), .C(n3609), .D(N7657), .Z(n238) );
  CND2X1 U11494 ( .A(N5780), .B(n3691), .Z(n237) );
  CANR2X1 U11495 ( .A(mem_data1[622]), .B(n3898), .C(N8902), .D(n3652), .Z(
        n236) );
  CND3XL U11496 ( .A(n239), .B(n240), .C(n241), .Z(N9945) );
  CANR2X1 U11497 ( .A(N2697), .B(n3574), .C(n3609), .D(N7658), .Z(n241) );
  CND2X1 U11498 ( .A(N5779), .B(n3697), .Z(n240) );
  CANR2X1 U11499 ( .A(mem_data1[621]), .B(n3898), .C(N8901), .D(n3652), .Z(
        n239) );
  CND3XL U11500 ( .A(n242), .B(n243), .C(n244), .Z(N9944) );
  CANR2X1 U11501 ( .A(N2696), .B(n3573), .C(n3609), .D(N7659), .Z(n244) );
  CND2X1 U11502 ( .A(N5778), .B(n3687), .Z(n243) );
  CANR2X1 U11503 ( .A(mem_data1[620]), .B(n3898), .C(N8900), .D(n3652), .Z(
        n242) );
  CND3XL U11504 ( .A(n245), .B(n246), .C(n247), .Z(N9943) );
  CANR2X1 U11505 ( .A(N2695), .B(n3573), .C(n3609), .D(N7660), .Z(n247) );
  CND2X1 U11506 ( .A(N5777), .B(n3688), .Z(n246) );
  CANR2X1 U11507 ( .A(mem_data1[619]), .B(n3898), .C(N8899), .D(n3652), .Z(
        n245) );
  CND3XL U11508 ( .A(n248), .B(n249), .C(n250), .Z(N9942) );
  CANR2X1 U11509 ( .A(N2694), .B(n3573), .C(n3609), .D(N7661), .Z(n250) );
  CND2X1 U11510 ( .A(N5776), .B(n3686), .Z(n249) );
  CANR2X1 U11511 ( .A(mem_data1[618]), .B(n3898), .C(N8898), .D(n3652), .Z(
        n248) );
  CND3XL U11512 ( .A(n251), .B(n252), .C(n253), .Z(N9941) );
  CANR2X1 U11513 ( .A(N2693), .B(n3573), .C(n3609), .D(N7662), .Z(n253) );
  CND2X1 U11514 ( .A(N5775), .B(n3696), .Z(n252) );
  CANR2X1 U11515 ( .A(mem_data1[617]), .B(n3898), .C(N8897), .D(n3654), .Z(
        n251) );
  CND3XL U11516 ( .A(n254), .B(n255), .C(n256), .Z(N9940) );
  CANR2X1 U11517 ( .A(N2692), .B(n3573), .C(n3609), .D(N7663), .Z(n256) );
  CND2X1 U11518 ( .A(N5774), .B(n3694), .Z(n255) );
  CANR2X1 U11519 ( .A(mem_data1[616]), .B(n3898), .C(N8896), .D(n3654), .Z(
        n254) );
  CND3XL U11520 ( .A(n257), .B(n258), .C(n259), .Z(N9939) );
  CANR2X1 U11521 ( .A(N2691), .B(n3573), .C(n3609), .D(N7664), .Z(n259) );
  CND2X1 U11522 ( .A(N5773), .B(n3695), .Z(n258) );
  CANR2X1 U11523 ( .A(mem_data1[615]), .B(n3898), .C(N8895), .D(n3654), .Z(
        n257) );
  CND3XL U11524 ( .A(n260), .B(n261), .C(n262), .Z(N9938) );
  CANR2X1 U11525 ( .A(N2690), .B(n3573), .C(n3609), .D(N7665), .Z(n262) );
  CND2X1 U11526 ( .A(N5772), .B(n3689), .Z(n261) );
  CANR2X1 U11527 ( .A(mem_data1[614]), .B(n3898), .C(N8894), .D(n3654), .Z(
        n260) );
  CND3XL U11528 ( .A(n263), .B(n264), .C(n265), .Z(N9937) );
  CANR2X1 U11529 ( .A(N2689), .B(n3573), .C(n3609), .D(N7666), .Z(n265) );
  CND2X1 U11530 ( .A(N5771), .B(n3698), .Z(n264) );
  CANR2X1 U11531 ( .A(mem_data1[613]), .B(n3898), .C(N8893), .D(n3654), .Z(
        n263) );
  CND3XL U11532 ( .A(n266), .B(n267), .C(n268), .Z(N9936) );
  CANR2X1 U11533 ( .A(N2688), .B(n3573), .C(n3609), .D(N7667), .Z(n268) );
  CND2X1 U11534 ( .A(N5770), .B(n3689), .Z(n267) );
  CANR2X1 U11535 ( .A(mem_data1[612]), .B(n3898), .C(N8892), .D(n3654), .Z(
        n266) );
  CND3XL U11536 ( .A(n269), .B(n270), .C(n271), .Z(N9935) );
  CANR2X1 U11537 ( .A(N2687), .B(n3573), .C(n3609), .D(N7668), .Z(n271) );
  CND2X1 U11538 ( .A(N5769), .B(n3696), .Z(n270) );
  CANR2X1 U11539 ( .A(mem_data1[611]), .B(n3898), .C(N8891), .D(n3654), .Z(
        n269) );
  CND3XL U11540 ( .A(n272), .B(n273), .C(n274), .Z(N9934) );
  CANR2X1 U11541 ( .A(N2686), .B(n3584), .C(n3609), .D(N7669), .Z(n274) );
  CND2X1 U11542 ( .A(N5768), .B(n3691), .Z(n273) );
  CANR2X1 U11543 ( .A(mem_data1[610]), .B(n3898), .C(N8890), .D(n3654), .Z(
        n272) );
  CND3XL U11544 ( .A(n275), .B(n276), .C(n277), .Z(N9933) );
  CANR2X1 U11545 ( .A(N2685), .B(n3584), .C(n3619), .D(N7670), .Z(n277) );
  CND2X1 U11546 ( .A(N5767), .B(n3687), .Z(n276) );
  CANR2X1 U11547 ( .A(mem_data1[609]), .B(n3898), .C(N8889), .D(n3654), .Z(
        n275) );
  CND3XL U11548 ( .A(n278), .B(n279), .C(n280), .Z(N9932) );
  CANR2X1 U11549 ( .A(N2684), .B(n3584), .C(n3619), .D(N7671), .Z(n280) );
  CND2X1 U11550 ( .A(N5766), .B(n3689), .Z(n279) );
  CANR2X1 U11551 ( .A(mem_data1[608]), .B(n3898), .C(N8888), .D(n3654), .Z(
        n278) );
  CND3XL U11552 ( .A(n281), .B(n282), .C(n283), .Z(N9931) );
  CANR2X1 U11553 ( .A(N2683), .B(n3584), .C(n3619), .D(N7672), .Z(n283) );
  CND2X1 U11554 ( .A(N5765), .B(n3691), .Z(n282) );
  CANR2X1 U11555 ( .A(mem_data1[607]), .B(n3898), .C(N8887), .D(n3654), .Z(
        n281) );
  CND3XL U11556 ( .A(n284), .B(n285), .C(n286), .Z(N9930) );
  CANR2X1 U11557 ( .A(N2682), .B(n3584), .C(n3619), .D(N7673), .Z(n286) );
  CND2X1 U11558 ( .A(N5764), .B(n3683), .Z(n285) );
  CANR2X1 U11559 ( .A(mem_data1[606]), .B(n3898), .C(N8886), .D(n3654), .Z(
        n284) );
  CND3XL U11560 ( .A(n287), .B(n288), .C(n289), .Z(N9929) );
  CANR2X1 U11561 ( .A(N2681), .B(n3584), .C(n3619), .D(N7674), .Z(n289) );
  CND2X1 U11562 ( .A(N5763), .B(n3688), .Z(n288) );
  CANR2X1 U11563 ( .A(mem_data1[605]), .B(n3898), .C(N8885), .D(n3654), .Z(
        n287) );
  CND3XL U11564 ( .A(n290), .B(n291), .C(n292), .Z(N9928) );
  CANR2X1 U11565 ( .A(N2680), .B(n3584), .C(n3619), .D(N7675), .Z(n292) );
  CND2X1 U11566 ( .A(N5762), .B(n3688), .Z(n291) );
  CANR2X1 U11567 ( .A(mem_data1[604]), .B(n3898), .C(N8884), .D(n3654), .Z(
        n290) );
  CND3XL U11568 ( .A(n293), .B(n294), .C(n295), .Z(N9927) );
  CANR2X1 U11569 ( .A(N2679), .B(n3584), .C(n3619), .D(N7676), .Z(n295) );
  CND2X1 U11570 ( .A(N5761), .B(n3688), .Z(n294) );
  CANR2X1 U11571 ( .A(mem_data1[603]), .B(n3898), .C(N8883), .D(n3654), .Z(
        n293) );
  CND3XL U11572 ( .A(n296), .B(n297), .C(n298), .Z(N9926) );
  CANR2X1 U11573 ( .A(N2678), .B(n3583), .C(n3619), .D(N7677), .Z(n298) );
  CND2X1 U11574 ( .A(N5760), .B(n3688), .Z(n297) );
  CANR2X1 U11575 ( .A(mem_data1[602]), .B(n3898), .C(N8882), .D(n3653), .Z(
        n296) );
  CND3XL U11576 ( .A(n299), .B(n300), .C(n301), .Z(N9925) );
  CANR2X1 U11577 ( .A(N2677), .B(n3583), .C(n3619), .D(N7678), .Z(n301) );
  CND2X1 U11578 ( .A(N5759), .B(n3688), .Z(n300) );
  CANR2X1 U11579 ( .A(mem_data1[601]), .B(n3898), .C(N8881), .D(n3653), .Z(
        n299) );
  CND3XL U11580 ( .A(n302), .B(n303), .C(n304), .Z(N9924) );
  CANR2X1 U11581 ( .A(N2676), .B(n3583), .C(n3619), .D(N7679), .Z(n304) );
  CND2X1 U11582 ( .A(N5758), .B(n3688), .Z(n303) );
  CANR2X1 U11583 ( .A(mem_data1[600]), .B(n3898), .C(N8880), .D(n3653), .Z(
        n302) );
  CND3XL U11584 ( .A(n305), .B(n306), .C(n307), .Z(N9923) );
  CANR2X1 U11585 ( .A(N2675), .B(n3583), .C(n3618), .D(N7680), .Z(n307) );
  CND2X1 U11586 ( .A(N5757), .B(n3688), .Z(n306) );
  CANR2X1 U11587 ( .A(mem_data1[599]), .B(n3898), .C(N8879), .D(n3653), .Z(
        n305) );
  CND3XL U11588 ( .A(n308), .B(n309), .C(n310), .Z(N9922) );
  CANR2X1 U11589 ( .A(N2674), .B(n3583), .C(n3618), .D(N7681), .Z(n310) );
  CND2X1 U11590 ( .A(N5756), .B(n3688), .Z(n309) );
  CANR2X1 U11591 ( .A(mem_data1[598]), .B(n3898), .C(N8878), .D(n3653), .Z(
        n308) );
  CND3XL U11592 ( .A(n311), .B(n312), .C(n313), .Z(N9921) );
  CANR2X1 U11593 ( .A(N2673), .B(n3583), .C(n3618), .D(N7682), .Z(n313) );
  CND2X1 U11594 ( .A(N5755), .B(n3688), .Z(n312) );
  CANR2X1 U11595 ( .A(mem_data1[597]), .B(n3898), .C(N8877), .D(n3653), .Z(
        n311) );
  CND3XL U11596 ( .A(n314), .B(n315), .C(n316), .Z(N9920) );
  CANR2X1 U11597 ( .A(N2672), .B(n3583), .C(n3618), .D(N7683), .Z(n316) );
  CND2X1 U11598 ( .A(N5754), .B(n3688), .Z(n315) );
  CANR2X1 U11599 ( .A(mem_data1[596]), .B(n3898), .C(N8876), .D(n3653), .Z(
        n314) );
  CND3XL U11600 ( .A(n317), .B(n318), .C(n319), .Z(N9919) );
  CANR2X1 U11601 ( .A(N2671), .B(n3583), .C(n3618), .D(N7684), .Z(n319) );
  CND2X1 U11602 ( .A(N5753), .B(n3696), .Z(n318) );
  CANR2X1 U11603 ( .A(mem_data1[595]), .B(n3898), .C(N8875), .D(n3655), .Z(
        n317) );
  CND3XL U11604 ( .A(n320), .B(n321), .C(n322), .Z(N9918) );
  CANR2X1 U11605 ( .A(N2670), .B(n3583), .C(n3618), .D(N7685), .Z(n322) );
  CND2X1 U11606 ( .A(N5752), .B(n3695), .Z(n321) );
  CANR2X1 U11607 ( .A(mem_data1[594]), .B(n3898), .C(N8874), .D(n3655), .Z(
        n320) );
  CND3XL U11608 ( .A(n323), .B(n324), .C(n325), .Z(N9917) );
  CANR2X1 U11609 ( .A(N2669), .B(n3583), .C(n3618), .D(N7686), .Z(n325) );
  CND2X1 U11610 ( .A(N5751), .B(n3687), .Z(n324) );
  CANR2X1 U11611 ( .A(mem_data1[593]), .B(n3898), .C(N8873), .D(n3655), .Z(
        n323) );
  CND3XL U11612 ( .A(n326), .B(n327), .C(n328), .Z(N9916) );
  CANR2X1 U11613 ( .A(N2668), .B(n3583), .C(n3618), .D(N7687), .Z(n328) );
  CND2X1 U11614 ( .A(N5750), .B(n3684), .Z(n327) );
  CANR2X1 U11615 ( .A(mem_data1[592]), .B(n3898), .C(N8872), .D(n3655), .Z(
        n326) );
  CND3XL U11616 ( .A(n329), .B(n330), .C(n331), .Z(N9915) );
  CANR2X1 U11617 ( .A(N2667), .B(n3583), .C(n3618), .D(N7688), .Z(n331) );
  CND2X1 U11618 ( .A(N5749), .B(n3693), .Z(n330) );
  CANR2X1 U11619 ( .A(mem_data1[591]), .B(n3898), .C(N8871), .D(n3655), .Z(
        n329) );
  CND3XL U11620 ( .A(n332), .B(n333), .C(n334), .Z(N9914) );
  CANR2X1 U11621 ( .A(N2666), .B(n3583), .C(n3618), .D(N7689), .Z(n334) );
  CND2X1 U11622 ( .A(N5748), .B(n3697), .Z(n333) );
  CANR2X1 U11623 ( .A(mem_data1[590]), .B(n3898), .C(N8870), .D(n3655), .Z(
        n332) );
  CND3XL U11624 ( .A(n335), .B(n336), .C(n337), .Z(N9913) );
  CANR2X1 U11625 ( .A(N2665), .B(n3583), .C(n3618), .D(N7690), .Z(n337) );
  CND2X1 U11626 ( .A(N5747), .B(n3697), .Z(n336) );
  CANR2X1 U11627 ( .A(mem_data1[589]), .B(n3898), .C(N8869), .D(n3655), .Z(
        n335) );
  CND3XL U11628 ( .A(n338), .B(n339), .C(n340), .Z(N9912) );
  CANR2X1 U11629 ( .A(N2664), .B(n3583), .C(n3618), .D(N7691), .Z(n340) );
  CND2X1 U11630 ( .A(N5746), .B(n3693), .Z(n339) );
  CANR2X1 U11631 ( .A(mem_data1[588]), .B(n3898), .C(N8868), .D(n3655), .Z(
        n338) );
  CND3XL U11632 ( .A(n341), .B(n342), .C(n343), .Z(N9911) );
  CANR2X1 U11633 ( .A(N2663), .B(n3583), .C(n3618), .D(N7692), .Z(n343) );
  CND2X1 U11634 ( .A(N5745), .B(n3683), .Z(n342) );
  CANR2X1 U11635 ( .A(mem_data1[587]), .B(n3898), .C(N8867), .D(n3655), .Z(
        n341) );
  CND3XL U11636 ( .A(n344), .B(n345), .C(n346), .Z(N9910) );
  CANR2X1 U11637 ( .A(N2662), .B(n3585), .C(n3618), .D(N7693), .Z(n346) );
  CND2X1 U11638 ( .A(N5744), .B(n3697), .Z(n345) );
  CANR2X1 U11639 ( .A(mem_data1[586]), .B(n3898), .C(N8866), .D(n3655), .Z(
        n344) );
  CND3XL U11640 ( .A(n347), .B(n348), .C(n349), .Z(N9909) );
  CANR2X1 U11641 ( .A(N2661), .B(n3585), .C(n3618), .D(N7694), .Z(n349) );
  CND2X1 U11642 ( .A(N5743), .B(n3683), .Z(n348) );
  CANR2X1 U11643 ( .A(mem_data1[585]), .B(n3898), .C(N8865), .D(n3655), .Z(
        n347) );
  CND3XL U11644 ( .A(n350), .B(n351), .C(n352), .Z(N9908) );
  CANR2X1 U11645 ( .A(N2660), .B(n3585), .C(n3618), .D(N7695), .Z(n352) );
  CND2X1 U11646 ( .A(N5742), .B(n3698), .Z(n351) );
  CANR2X1 U11647 ( .A(mem_data1[584]), .B(n3898), .C(N8864), .D(n3655), .Z(
        n350) );
  CND3XL U11648 ( .A(n353), .B(n354), .C(n355), .Z(N9907) );
  CANR2X1 U11649 ( .A(N2659), .B(n3585), .C(n3618), .D(N7696), .Z(n355) );
  CND2X1 U11650 ( .A(N5741), .B(n3698), .Z(n354) );
  CANR2X1 U11651 ( .A(mem_data1[583]), .B(n3898), .C(N8863), .D(n3655), .Z(
        n353) );
  CND3XL U11652 ( .A(n356), .B(n357), .C(n358), .Z(N9906) );
  CANR2X1 U11653 ( .A(N2658), .B(n3585), .C(n3620), .D(N7697), .Z(n358) );
  CND2X1 U11654 ( .A(N5740), .B(n3690), .Z(n357) );
  CANR2X1 U11655 ( .A(mem_data1[582]), .B(n3898), .C(N8862), .D(n3655), .Z(
        n356) );
  CND3XL U11656 ( .A(n359), .B(n360), .C(n361), .Z(N9905) );
  CANR2X1 U11657 ( .A(N2657), .B(n3585), .C(n3620), .D(N7698), .Z(n361) );
  CND2X1 U11658 ( .A(N5739), .B(n3696), .Z(n360) );
  CANR2X1 U11659 ( .A(mem_data1[581]), .B(n3898), .C(N8861), .D(n3655), .Z(
        n359) );
  CND3XL U11660 ( .A(n362), .B(n363), .C(n364), .Z(N9904) );
  CANR2X1 U11661 ( .A(N2656), .B(n3585), .C(n3620), .D(N7699), .Z(n364) );
  CND2X1 U11662 ( .A(N5738), .B(n3694), .Z(n363) );
  CANR2X1 U11663 ( .A(mem_data1[580]), .B(n3898), .C(N8860), .D(n3654), .Z(
        n362) );
  CND3XL U11664 ( .A(n365), .B(n366), .C(n367), .Z(N9903) );
  CANR2X1 U11665 ( .A(N2655), .B(n3585), .C(n3620), .D(N7700), .Z(n367) );
  CND2X1 U11666 ( .A(N5737), .B(n3695), .Z(n366) );
  CANR2X1 U11667 ( .A(mem_data1[579]), .B(n3898), .C(N8859), .D(n3654), .Z(
        n365) );
  CND3XL U11668 ( .A(n368), .B(n369), .C(n370), .Z(N9902) );
  CANR2X1 U11669 ( .A(N2654), .B(n3585), .C(n3620), .D(N7701), .Z(n370) );
  CND2X1 U11670 ( .A(N5736), .B(n3684), .Z(n369) );
  CANR2X1 U11671 ( .A(mem_data1[578]), .B(n3898), .C(N8858), .D(n3654), .Z(
        n368) );
  CND3XL U11672 ( .A(n371), .B(n372), .C(n373), .Z(N9901) );
  CANR2X1 U11673 ( .A(N2653), .B(n3584), .C(n3620), .D(N7702), .Z(n373) );
  CND2X1 U11674 ( .A(N5735), .B(n3690), .Z(n372) );
  CANR2X1 U11675 ( .A(mem_data1[577]), .B(n3898), .C(N8857), .D(n3654), .Z(
        n371) );
  CND3XL U11676 ( .A(n374), .B(n375), .C(n376), .Z(N9900) );
  CANR2X1 U11677 ( .A(N2652), .B(n3584), .C(n3620), .D(N7703), .Z(n376) );
  CND2X1 U11678 ( .A(N5734), .B(n3689), .Z(n375) );
  CANR2X1 U11679 ( .A(mem_data1[576]), .B(n3898), .C(N8856), .D(n3654), .Z(
        n374) );
  CND3XL U11680 ( .A(n377), .B(n378), .C(n379), .Z(N9899) );
  CANR2X1 U11681 ( .A(N2651), .B(n3584), .C(n3620), .D(N7704), .Z(n379) );
  CND2X1 U11682 ( .A(N5733), .B(n3694), .Z(n378) );
  CANR2X1 U11683 ( .A(mem_data1[575]), .B(n3898), .C(N8855), .D(n3654), .Z(
        n377) );
  CND3XL U11684 ( .A(n380), .B(n381), .C(n382), .Z(N9898) );
  CANR2X1 U11685 ( .A(N2650), .B(n3584), .C(n3620), .D(N7705), .Z(n382) );
  CND2X1 U11686 ( .A(N5732), .B(n3697), .Z(n381) );
  CANR2X1 U11687 ( .A(mem_data1[574]), .B(n3898), .C(N8854), .D(n3654), .Z(
        n380) );
  CND3XL U11688 ( .A(n383), .B(n384), .C(n385), .Z(N9897) );
  CANR2X1 U11689 ( .A(N2649), .B(n3584), .C(n3620), .D(N7706), .Z(n385) );
  CND2X1 U11690 ( .A(N5731), .B(n3690), .Z(n384) );
  CANR2X1 U11691 ( .A(mem_data1[573]), .B(n3898), .C(N8853), .D(n3656), .Z(
        n383) );
  CND3XL U11692 ( .A(n386), .B(n387), .C(n388), .Z(N9896) );
  CANR2X1 U11693 ( .A(N2648), .B(n3584), .C(n3619), .D(N7707), .Z(n388) );
  CND2X1 U11694 ( .A(N5730), .B(n3690), .Z(n387) );
  CANR2X1 U11695 ( .A(mem_data1[572]), .B(n3898), .C(N8852), .D(n3656), .Z(
        n386) );
  CND3XL U11696 ( .A(n389), .B(n390), .C(n391), .Z(N9895) );
  CANR2X1 U11697 ( .A(N2647), .B(n3584), .C(n3619), .D(N7708), .Z(n391) );
  CND2X1 U11698 ( .A(N5729), .B(n3695), .Z(n390) );
  CANR2X1 U11699 ( .A(mem_data1[571]), .B(n3898), .C(N8851), .D(n3656), .Z(
        n389) );
  CND3XL U11700 ( .A(n392), .B(n393), .C(n394), .Z(N9894) );
  CANR2X1 U11701 ( .A(N2646), .B(n3584), .C(n3619), .D(N7709), .Z(n394) );
  CND2X1 U11702 ( .A(N5728), .B(n3689), .Z(n393) );
  CANR2X1 U11703 ( .A(mem_data1[570]), .B(n3898), .C(N8850), .D(n3656), .Z(
        n392) );
  CND3XL U11704 ( .A(n395), .B(n396), .C(n397), .Z(N9893) );
  CANR2X1 U11705 ( .A(N2645), .B(n3584), .C(n3619), .D(N7710), .Z(n397) );
  CND2X1 U11706 ( .A(N5727), .B(n3686), .Z(n396) );
  CANR2X1 U11707 ( .A(mem_data1[569]), .B(n3898), .C(N8849), .D(n3656), .Z(
        n395) );
  CND3XL U11708 ( .A(n398), .B(n399), .C(n400), .Z(N9892) );
  CANR2X1 U11709 ( .A(N2644), .B(n3584), .C(n3619), .D(N7711), .Z(n400) );
  CND2X1 U11710 ( .A(N5726), .B(n3689), .Z(n399) );
  CANR2X1 U11711 ( .A(mem_data1[568]), .B(n3898), .C(N8848), .D(n3656), .Z(
        n398) );
  CND3XL U11712 ( .A(n401), .B(n402), .C(n403), .Z(N9891) );
  CANR2X1 U11713 ( .A(N2643), .B(n3584), .C(n3619), .D(N7712), .Z(n403) );
  CND2X1 U11714 ( .A(N5725), .B(n3685), .Z(n402) );
  CANR2X1 U11715 ( .A(mem_data1[567]), .B(n3898), .C(N8847), .D(n3656), .Z(
        n401) );
  CND3XL U11716 ( .A(n404), .B(n405), .C(n406), .Z(N9890) );
  CANR2X1 U11717 ( .A(N2642), .B(n3584), .C(n3619), .D(N7713), .Z(n406) );
  CND2X1 U11718 ( .A(N5724), .B(n3693), .Z(n405) );
  CANR2X1 U11719 ( .A(mem_data1[566]), .B(n3898), .C(N8846), .D(n3656), .Z(
        n404) );
  CND3XL U11720 ( .A(n407), .B(n408), .C(n409), .Z(N9889) );
  CANR2X1 U11721 ( .A(N2641), .B(n3584), .C(n3619), .D(N7714), .Z(n409) );
  CND2X1 U11722 ( .A(N5723), .B(n3687), .Z(n408) );
  CANR2X1 U11723 ( .A(mem_data1[565]), .B(n3898), .C(N8845), .D(n3656), .Z(
        n407) );
  CND3XL U11724 ( .A(n410), .B(n411), .C(n412), .Z(N9888) );
  CANR2X1 U11725 ( .A(N2640), .B(n3584), .C(n3619), .D(N7715), .Z(n412) );
  CND2X1 U11726 ( .A(N5722), .B(n3689), .Z(n411) );
  CANR2X1 U11727 ( .A(mem_data1[564]), .B(n3898), .C(N8844), .D(n3656), .Z(
        n410) );
  CND3XL U11728 ( .A(n413), .B(n414), .C(n415), .Z(N9887) );
  CANR2X1 U11729 ( .A(N2639), .B(n3584), .C(n3619), .D(N7716), .Z(n415) );
  CND2X1 U11730 ( .A(N5721), .B(n3683), .Z(n414) );
  CANR2X1 U11731 ( .A(mem_data1[563]), .B(n3898), .C(N8843), .D(n3656), .Z(
        n413) );
  CND3XL U11732 ( .A(n416), .B(n417), .C(n418), .Z(N9886) );
  CANR2X1 U11733 ( .A(N2638), .B(n3584), .C(n3619), .D(N7717), .Z(n418) );
  CND2X1 U11734 ( .A(N5720), .B(n3691), .Z(n417) );
  CANR2X1 U11735 ( .A(mem_data1[562]), .B(n3898), .C(N8842), .D(n3656), .Z(
        n416) );
  CND3XL U11736 ( .A(n419), .B(n420), .C(n421), .Z(N9885) );
  CANR2X1 U11737 ( .A(N2637), .B(n3586), .C(n3619), .D(N7718), .Z(n421) );
  CND2X1 U11738 ( .A(N5719), .B(n3684), .Z(n420) );
  CANR2X1 U11739 ( .A(mem_data1[561]), .B(n3898), .C(N8841), .D(n3656), .Z(
        n419) );
  CND3XL U11740 ( .A(n422), .B(n423), .C(n424), .Z(N9884) );
  CANR2X1 U11741 ( .A(N2636), .B(n3586), .C(n3619), .D(N7719), .Z(n424) );
  CND2X1 U11742 ( .A(N5718), .B(n3687), .Z(n423) );
  CANR2X1 U11743 ( .A(mem_data1[560]), .B(n3898), .C(N8840), .D(n3656), .Z(
        n422) );
  CND3XL U11744 ( .A(n425), .B(n426), .C(n427), .Z(N9883) );
  CANR2X1 U11745 ( .A(N2635), .B(n3586), .C(n3619), .D(N7720), .Z(n427) );
  CND2X1 U11746 ( .A(N5717), .B(n3697), .Z(n426) );
  CANR2X1 U11747 ( .A(mem_data1[559]), .B(n3898), .C(N8839), .D(n3656), .Z(
        n425) );
  CND3XL U11748 ( .A(n428), .B(n429), .C(n430), .Z(N9882) );
  CANR2X1 U11749 ( .A(N2634), .B(n3586), .C(n3619), .D(N7721), .Z(n430) );
  CND2X1 U11750 ( .A(N5716), .B(n3686), .Z(n429) );
  CANR2X1 U11751 ( .A(mem_data1[558]), .B(n3898), .C(N8838), .D(n3656), .Z(
        n428) );
  CND3XL U11752 ( .A(n431), .B(n432), .C(n433), .Z(N9881) );
  CANR2X1 U11753 ( .A(N2633), .B(n3586), .C(n3619), .D(N7722), .Z(n433) );
  CND2X1 U11754 ( .A(N5715), .B(n3693), .Z(n432) );
  CANR2X1 U11755 ( .A(mem_data1[557]), .B(n3898), .C(N8837), .D(n3655), .Z(
        n431) );
  CND3XL U11756 ( .A(n434), .B(n435), .C(n436), .Z(N9880) );
  CANR2X1 U11757 ( .A(N2632), .B(n3586), .C(n3619), .D(N7723), .Z(n436) );
  CND2X1 U11758 ( .A(N5714), .B(n3697), .Z(n435) );
  CANR2X1 U11759 ( .A(mem_data1[556]), .B(n3898), .C(N8836), .D(n3655), .Z(
        n434) );
  CND3XL U11760 ( .A(n437), .B(n438), .C(n439), .Z(N9879) );
  CANR2X1 U11761 ( .A(N2631), .B(n3586), .C(n3621), .D(N7724), .Z(n439) );
  CND2X1 U11762 ( .A(N5713), .B(n3697), .Z(n438) );
  CANR2X1 U11763 ( .A(mem_data1[555]), .B(n3898), .C(N8835), .D(n3655), .Z(
        n437) );
  CND3XL U11764 ( .A(n440), .B(n441), .C(n442), .Z(N9878) );
  CANR2X1 U11765 ( .A(N2630), .B(n3587), .C(n3621), .D(N7725), .Z(n442) );
  CND2X1 U11766 ( .A(N5712), .B(n3695), .Z(n441) );
  CANR2X1 U11767 ( .A(mem_data1[554]), .B(n3898), .C(N8834), .D(n3655), .Z(
        n440) );
  CND3XL U11768 ( .A(n443), .B(n444), .C(n445), .Z(N9877) );
  CANR2X1 U11769 ( .A(N2629), .B(n3585), .C(n3621), .D(N7726), .Z(n445) );
  CND2X1 U11770 ( .A(N5711), .B(n3689), .Z(n444) );
  CANR2X1 U11771 ( .A(mem_data1[553]), .B(n3898), .C(N8833), .D(n3655), .Z(
        n443) );
  CND3XL U11772 ( .A(n446), .B(n447), .C(n448), .Z(N9876) );
  CANR2X1 U11773 ( .A(N2628), .B(n3585), .C(n3621), .D(N7727), .Z(n448) );
  CND2X1 U11774 ( .A(N5710), .B(n3683), .Z(n447) );
  CANR2X1 U11775 ( .A(mem_data1[552]), .B(n3898), .C(N8832), .D(n3655), .Z(
        n446) );
  CND3XL U11776 ( .A(n449), .B(n450), .C(n451), .Z(N9875) );
  CANR2X1 U11777 ( .A(N2627), .B(n3585), .C(n3621), .D(N7728), .Z(n451) );
  CND2X1 U11778 ( .A(N5709), .B(n3685), .Z(n450) );
  CANR2X1 U11779 ( .A(mem_data1[551]), .B(n3898), .C(N8831), .D(n3657), .Z(
        n449) );
  CND3XL U11780 ( .A(n452), .B(n453), .C(n454), .Z(N9874) );
  CANR2X1 U11781 ( .A(N2626), .B(n3585), .C(n3620), .D(N7729), .Z(n454) );
  CND2X1 U11782 ( .A(N5708), .B(n3685), .Z(n453) );
  CANR2X1 U11783 ( .A(mem_data1[550]), .B(n3898), .C(N8830), .D(n3657), .Z(
        n452) );
  CND3XL U11784 ( .A(n455), .B(n456), .C(n457), .Z(N9873) );
  CANR2X1 U11785 ( .A(N2625), .B(n3585), .C(n3620), .D(N7730), .Z(n457) );
  CND2X1 U11786 ( .A(N5707), .B(n3685), .Z(n456) );
  CANR2X1 U11787 ( .A(mem_data1[549]), .B(n3898), .C(N8829), .D(n3657), .Z(
        n455) );
  CND3XL U11788 ( .A(n458), .B(n459), .C(n460), .Z(N9872) );
  CANR2X1 U11789 ( .A(N2624), .B(n3585), .C(n3620), .D(N7731), .Z(n460) );
  CND2X1 U11790 ( .A(N5706), .B(n3685), .Z(n459) );
  CANR2X1 U11791 ( .A(mem_data1[548]), .B(n3898), .C(N8828), .D(n3657), .Z(
        n458) );
  CND3XL U11792 ( .A(n461), .B(n462), .C(n463), .Z(N9871) );
  CANR2X1 U11793 ( .A(N2623), .B(n3584), .C(n3620), .D(N7732), .Z(n463) );
  CND2X1 U11794 ( .A(N5705), .B(n3685), .Z(n462) );
  CANR2X1 U11795 ( .A(mem_data1[547]), .B(n3898), .C(N8827), .D(n3657), .Z(
        n461) );
  CND3XL U11796 ( .A(n464), .B(n465), .C(n466), .Z(N9870) );
  CANR2X1 U11797 ( .A(N2622), .B(n3578), .C(n3609), .D(N7733), .Z(n466) );
  CND2X1 U11798 ( .A(N5704), .B(n3685), .Z(n465) );
  CANR2X1 U11799 ( .A(mem_data1[546]), .B(n3898), .C(N8826), .D(n3657), .Z(
        n464) );
  CND3XL U11800 ( .A(n467), .B(n468), .C(n469), .Z(N9869) );
  CANR2X1 U11801 ( .A(N2621), .B(n3578), .C(n3612), .D(N7734), .Z(n469) );
  CND2X1 U11802 ( .A(N5703), .B(n3685), .Z(n468) );
  CANR2X1 U11803 ( .A(mem_data1[545]), .B(n3898), .C(N8825), .D(n3657), .Z(
        n467) );
  CND3XL U11804 ( .A(n470), .B(n471), .C(n472), .Z(N9868) );
  CANR2X1 U11805 ( .A(N2620), .B(n3577), .C(n3612), .D(N7735), .Z(n472) );
  CND2X1 U11806 ( .A(N5702), .B(n3685), .Z(n471) );
  CANR2X1 U11807 ( .A(mem_data1[544]), .B(n3898), .C(N8824), .D(n3657), .Z(
        n470) );
  CND3XL U11808 ( .A(n473), .B(n474), .C(n475), .Z(N9867) );
  CANR2X1 U11809 ( .A(N2619), .B(n3577), .C(n3612), .D(N7736), .Z(n475) );
  CND2X1 U11810 ( .A(N5701), .B(n3685), .Z(n474) );
  CANR2X1 U11811 ( .A(mem_data1[543]), .B(n3898), .C(N8823), .D(n3657), .Z(
        n473) );
  CND3XL U11812 ( .A(n476), .B(n477), .C(n478), .Z(N9866) );
  CANR2X1 U11813 ( .A(N2618), .B(n3577), .C(n3612), .D(N7737), .Z(n478) );
  CND2X1 U11814 ( .A(N5700), .B(n3685), .Z(n477) );
  CANR2X1 U11815 ( .A(mem_data1[542]), .B(n3898), .C(N8822), .D(n3657), .Z(
        n476) );
  CND3XL U11816 ( .A(n479), .B(n480), .C(n481), .Z(N9865) );
  CANR2X1 U11817 ( .A(N2617), .B(n3577), .C(n3612), .D(N7738), .Z(n481) );
  CND2X1 U11818 ( .A(N5699), .B(n3685), .Z(n480) );
  CANR2X1 U11819 ( .A(mem_data1[541]), .B(n3898), .C(N8821), .D(n3657), .Z(
        n479) );
  CND3XL U11820 ( .A(n482), .B(n483), .C(n484), .Z(N9864) );
  CANR2X1 U11821 ( .A(N2616), .B(n3577), .C(n3612), .D(N7739), .Z(n484) );
  CND2X1 U11822 ( .A(N5698), .B(n3685), .Z(n483) );
  CANR2X1 U11823 ( .A(mem_data1[540]), .B(n3898), .C(N8820), .D(n3657), .Z(
        n482) );
  CND3XL U11824 ( .A(n485), .B(n486), .C(n487), .Z(N9863) );
  CANR2X1 U11825 ( .A(N2615), .B(n3577), .C(n3608), .D(N7740), .Z(n487) );
  CND2X1 U11826 ( .A(N5697), .B(n3685), .Z(n486) );
  CANR2X1 U11827 ( .A(mem_data1[539]), .B(n3898), .C(N8819), .D(n3657), .Z(
        n485) );
  CND3XL U11828 ( .A(n488), .B(n489), .C(n490), .Z(N9862) );
  CANR2X1 U11829 ( .A(N2614), .B(n3577), .C(n3614), .D(N7741), .Z(n490) );
  CND2X1 U11830 ( .A(N5696), .B(n3685), .Z(n489) );
  CANR2X1 U11831 ( .A(mem_data1[538]), .B(n3898), .C(N8818), .D(n3657), .Z(
        n488) );
  CND3XL U11832 ( .A(n491), .B(n492), .C(n493), .Z(N9861) );
  CANR2X1 U11833 ( .A(N2613), .B(n3577), .C(n3614), .D(N7742), .Z(n493) );
  CND2X1 U11834 ( .A(N5695), .B(n3685), .Z(n492) );
  CANR2X1 U11835 ( .A(mem_data1[537]), .B(n3898), .C(N8817), .D(n3657), .Z(
        n491) );
  CND3XL U11836 ( .A(n494), .B(n495), .C(n496), .Z(N9860) );
  CANR2X1 U11837 ( .A(N2612), .B(n3577), .C(n3614), .D(N7743), .Z(n496) );
  CND2X1 U11838 ( .A(N5694), .B(n3685), .Z(n495) );
  CANR2X1 U11839 ( .A(mem_data1[536]), .B(n3898), .C(N8816), .D(n3657), .Z(
        n494) );
  CND3XL U11840 ( .A(n497), .B(n498), .C(n499), .Z(N9859) );
  CANR2X1 U11841 ( .A(N2611), .B(n3577), .C(n3614), .D(N7744), .Z(n499) );
  CND2X1 U11842 ( .A(N5693), .B(n3685), .Z(n498) );
  CANR2X1 U11843 ( .A(mem_data1[535]), .B(n3898), .C(N8815), .D(n3656), .Z(
        n497) );
  CND3XL U11844 ( .A(n500), .B(n501), .C(n502), .Z(N9858) );
  CANR2X1 U11845 ( .A(N2610), .B(n3577), .C(n3614), .D(N7745), .Z(n502) );
  CND2X1 U11846 ( .A(N5692), .B(n3685), .Z(n501) );
  CANR2X1 U11847 ( .A(mem_data1[534]), .B(n3898), .C(N8814), .D(n3656), .Z(
        n500) );
  CND3XL U11848 ( .A(n503), .B(n504), .C(n505), .Z(N9857) );
  CANR2X1 U11849 ( .A(N2609), .B(n3577), .C(n3613), .D(N7746), .Z(n505) );
  CND2X1 U11850 ( .A(N5691), .B(n3685), .Z(n504) );
  CANR2X1 U11851 ( .A(mem_data1[533]), .B(n3898), .C(N8813), .D(n3656), .Z(
        n503) );
  CND3XL U11852 ( .A(n506), .B(n507), .C(n508), .Z(N9856) );
  CANR2X1 U11853 ( .A(N2608), .B(n3577), .C(n3613), .D(N7747), .Z(n508) );
  CND2X1 U11854 ( .A(N5690), .B(n3685), .Z(n507) );
  CANR2X1 U11855 ( .A(mem_data1[532]), .B(n3898), .C(N8812), .D(n3656), .Z(
        n506) );
  CND3XL U11856 ( .A(n509), .B(n510), .C(n511), .Z(N9855) );
  CANR2X1 U11857 ( .A(N2607), .B(n3577), .C(n3613), .D(N7748), .Z(n511) );
  CND2X1 U11858 ( .A(N5689), .B(n3693), .Z(n510) );
  CANR2X1 U11859 ( .A(mem_data1[531]), .B(n3898), .C(N8811), .D(n3656), .Z(
        n509) );
  CND3XL U11860 ( .A(n512), .B(n513), .C(n514), .Z(N9854) );
  CANR2X1 U11861 ( .A(N2606), .B(n3577), .C(n3613), .D(N7749), .Z(n514) );
  CND2X1 U11862 ( .A(N5688), .B(n3684), .Z(n513) );
  CANR2X1 U11863 ( .A(mem_data1[530]), .B(n3898), .C(N8810), .D(n3656), .Z(
        n512) );
  CND3XL U11864 ( .A(n515), .B(n516), .C(n517), .Z(N9853) );
  CANR2X1 U11865 ( .A(N2605), .B(n3577), .C(n3613), .D(N7750), .Z(n517) );
  CND2X1 U11866 ( .A(N5687), .B(n3690), .Z(n516) );
  CANR2X1 U11867 ( .A(mem_data1[529]), .B(n3898), .C(N8809), .D(n3658), .Z(
        n515) );
  CND3XL U11868 ( .A(n518), .B(n519), .C(n520), .Z(N9852) );
  CANR2X1 U11869 ( .A(N2604), .B(n3577), .C(n3613), .D(N7751), .Z(n520) );
  CND2X1 U11870 ( .A(N5686), .B(n3696), .Z(n519) );
  CANR2X1 U11871 ( .A(mem_data1[528]), .B(n3898), .C(N8808), .D(n3658), .Z(
        n518) );
  CND3XL U11872 ( .A(n521), .B(n522), .C(n523), .Z(N9851) );
  CANR2X1 U11873 ( .A(N2603), .B(n3570), .C(n3613), .D(N7752), .Z(n523) );
  CND2X1 U11874 ( .A(N5685), .B(n3694), .Z(n522) );
  CANR2X1 U11875 ( .A(mem_data1[527]), .B(n3898), .C(N8807), .D(n3658), .Z(
        n521) );
  CND3XL U11876 ( .A(n524), .B(n525), .C(n526), .Z(N9850) );
  CANR2X1 U11877 ( .A(N2602), .B(n3570), .C(n3613), .D(N7753), .Z(n526) );
  CND2X1 U11878 ( .A(N5684), .B(n3695), .Z(n525) );
  CANR2X1 U11879 ( .A(mem_data1[526]), .B(n3898), .C(N8806), .D(n3658), .Z(
        n524) );
  CND3XL U11880 ( .A(n527), .B(n528), .C(n529), .Z(N9849) );
  CANR2X1 U11881 ( .A(N2601), .B(n3570), .C(n3613), .D(N7754), .Z(n529) );
  CND2X1 U11882 ( .A(N5683), .B(n3697), .Z(n528) );
  CANR2X1 U11883 ( .A(mem_data1[525]), .B(n3898), .C(N8805), .D(n3658), .Z(
        n527) );
  CND3XL U11884 ( .A(n530), .B(n531), .C(n532), .Z(N9848) );
  CANR2X1 U11885 ( .A(N2600), .B(n3570), .C(n3613), .D(N7755), .Z(n532) );
  CND2X1 U11886 ( .A(N5682), .B(n3695), .Z(n531) );
  CANR2X1 U11887 ( .A(mem_data1[524]), .B(n3898), .C(N8804), .D(n3658), .Z(
        n530) );
  CND3XL U11888 ( .A(n533), .B(n534), .C(n535), .Z(N9847) );
  CANR2X1 U11889 ( .A(N2599), .B(n3570), .C(n3613), .D(N7756), .Z(n535) );
  CND2X1 U11890 ( .A(N5681), .B(n3689), .Z(n534) );
  CANR2X1 U11891 ( .A(mem_data1[523]), .B(n3898), .C(N8803), .D(n3658), .Z(
        n533) );
  CND3XL U11892 ( .A(n536), .B(n537), .C(n538), .Z(N9846) );
  CANR2X1 U11893 ( .A(N2598), .B(n3570), .C(n3613), .D(N7757), .Z(n538) );
  CND2X1 U11894 ( .A(N5680), .B(n3689), .Z(n537) );
  CANR2X1 U11895 ( .A(mem_data1[522]), .B(n3898), .C(N8802), .D(n3658), .Z(
        n536) );
  CND3XL U11896 ( .A(n539), .B(n540), .C(n541), .Z(N9845) );
  CANR2X1 U11897 ( .A(N2597), .B(n3570), .C(n3613), .D(N7758), .Z(n541) );
  CND2X1 U11898 ( .A(N5679), .B(n3690), .Z(n540) );
  CANR2X1 U11899 ( .A(mem_data1[521]), .B(n3898), .C(N8801), .D(n3658), .Z(
        n539) );
  CND3XL U11900 ( .A(n542), .B(n543), .C(n544), .Z(N9844) );
  CANR2X1 U11901 ( .A(N2596), .B(n3570), .C(n3613), .D(N7759), .Z(n544) );
  CND2X1 U11902 ( .A(N5678), .B(n3695), .Z(n543) );
  CANR2X1 U11903 ( .A(mem_data1[520]), .B(n3898), .C(N8800), .D(n3658), .Z(
        n542) );
  CND3XL U11904 ( .A(n545), .B(n546), .C(n547), .Z(N9843) );
  CANR2X1 U11905 ( .A(N2595), .B(n3570), .C(n3613), .D(N7760), .Z(n547) );
  CND2X1 U11906 ( .A(N5677), .B(n3698), .Z(n546) );
  CANR2X1 U11907 ( .A(mem_data1[519]), .B(n3898), .C(N8799), .D(n3658), .Z(
        n545) );
  CND3XL U11908 ( .A(n548), .B(n549), .C(n550), .Z(N9842) );
  CANR2X1 U11909 ( .A(N2594), .B(n3570), .C(n3613), .D(N7761), .Z(n550) );
  CND2X1 U11910 ( .A(N5676), .B(n3695), .Z(n549) );
  CANR2X1 U11911 ( .A(mem_data1[518]), .B(n3898), .C(N8798), .D(n3658), .Z(
        n548) );
  CND3XL U11912 ( .A(n551), .B(n552), .C(n553), .Z(N9841) );
  CANR2X1 U11913 ( .A(N2593), .B(n3572), .C(n3613), .D(N7762), .Z(n553) );
  CND2X1 U11914 ( .A(N5675), .B(n3684), .Z(n552) );
  CANR2X1 U11915 ( .A(mem_data1[517]), .B(n3898), .C(N8797), .D(n3658), .Z(
        n551) );
  CND3XL U11916 ( .A(n554), .B(n555), .C(n556), .Z(N9840) );
  CANR2X1 U11917 ( .A(N2592), .B(n3578), .C(n3613), .D(N7763), .Z(n556) );
  CND2X1 U11918 ( .A(N5674), .B(n3686), .Z(n555) );
  CANR2X1 U11919 ( .A(mem_data1[516]), .B(n3898), .C(N8796), .D(n3658), .Z(
        n554) );
  CND3XL U11920 ( .A(n557), .B(n558), .C(n559), .Z(N9839) );
  CANR2X1 U11921 ( .A(N2591), .B(n3578), .C(n3613), .D(N7764), .Z(n559) );
  CND2X1 U11922 ( .A(N5673), .B(n3697), .Z(n558) );
  CANR2X1 U11923 ( .A(mem_data1[515]), .B(n3898), .C(N8795), .D(n3658), .Z(
        n557) );
  CND3XL U11924 ( .A(n560), .B(n561), .C(n562), .Z(N9838) );
  CANR2X1 U11925 ( .A(N2590), .B(n3578), .C(n3613), .D(N7765), .Z(n562) );
  CND2X1 U11926 ( .A(N5672), .B(n3687), .Z(n561) );
  CANR2X1 U11927 ( .A(mem_data1[514]), .B(n3898), .C(N8794), .D(n3658), .Z(
        n560) );
  CND3XL U11928 ( .A(n563), .B(n564), .C(n565), .Z(N9837) );
  CANR2X1 U11929 ( .A(N2589), .B(n3578), .C(n3613), .D(N7766), .Z(n565) );
  CND2X1 U11930 ( .A(N5671), .B(n3691), .Z(n564) );
  CANR2X1 U11931 ( .A(mem_data1[513]), .B(n3898), .C(N8793), .D(n3657), .Z(
        n563) );
  CND3XL U11932 ( .A(n566), .B(n567), .C(n568), .Z(N9836) );
  CANR2X1 U11933 ( .A(N2588), .B(n3578), .C(n3606), .D(N7767), .Z(n568) );
  CND2X1 U11934 ( .A(N5670), .B(n3694), .Z(n567) );
  CANR2X1 U11935 ( .A(mem_data1[512]), .B(n3898), .C(N8792), .D(n3657), .Z(
        n566) );
  CND3XL U11936 ( .A(n569), .B(n570), .C(n571), .Z(N9835) );
  CANR2X1 U11937 ( .A(N2587), .B(n3578), .C(n3606), .D(N7768), .Z(n571) );
  CND2X1 U11938 ( .A(N5669), .B(n3690), .Z(n570) );
  CANR2X1 U11939 ( .A(mem_data1[511]), .B(n3898), .C(N8791), .D(n3657), .Z(
        n569) );
  CND3XL U11940 ( .A(n572), .B(n573), .C(n574), .Z(N9834) );
  CANR2X1 U11941 ( .A(N2586), .B(n3578), .C(n3606), .D(N7769), .Z(n574) );
  CND2X1 U11942 ( .A(N5668), .B(n3696), .Z(n573) );
  CANR2X1 U11943 ( .A(mem_data1[510]), .B(n3898), .C(N8790), .D(n3657), .Z(
        n572) );
  CND3XL U11944 ( .A(n575), .B(n576), .C(n577), .Z(N9833) );
  CANR2X1 U11945 ( .A(N2585), .B(n3578), .C(n3606), .D(N7770), .Z(n577) );
  CND2X1 U11946 ( .A(N5667), .B(n3685), .Z(n576) );
  CANR2X1 U11947 ( .A(mem_data1[509]), .B(n3898), .C(N8789), .D(n3657), .Z(
        n575) );
  CND3XL U11948 ( .A(n578), .B(n579), .C(n580), .Z(N9832) );
  CANR2X1 U11949 ( .A(N2584), .B(n3578), .C(n3606), .D(N7771), .Z(n580) );
  CND2X1 U11950 ( .A(N5666), .B(n3685), .Z(n579) );
  CANR2X1 U11951 ( .A(mem_data1[508]), .B(n3898), .C(N8788), .D(n3657), .Z(
        n578) );
  CND3XL U11952 ( .A(n581), .B(n582), .C(n583), .Z(N9831) );
  CANR2X1 U11953 ( .A(N2583), .B(n3578), .C(n3606), .D(N7772), .Z(n583) );
  CND2X1 U11954 ( .A(N5665), .B(n3686), .Z(n582) );
  CANR2X1 U11955 ( .A(mem_data1[507]), .B(n3898), .C(N8787), .D(n3659), .Z(
        n581) );
  CND3XL U11956 ( .A(n584), .B(n585), .C(n586), .Z(N9830) );
  CANR2X1 U11957 ( .A(N2582), .B(n3578), .C(n3606), .D(N7773), .Z(n586) );
  CND2X1 U11958 ( .A(N5664), .B(n3686), .Z(n585) );
  CANR2X1 U11959 ( .A(mem_data1[506]), .B(n3898), .C(N8786), .D(n3659), .Z(
        n584) );
  CND3XL U11960 ( .A(n587), .B(n588), .C(n589), .Z(N9829) );
  CANR2X1 U11961 ( .A(N2581), .B(n3578), .C(n3606), .D(N7774), .Z(n589) );
  CND2X1 U11962 ( .A(N5663), .B(n3686), .Z(n588) );
  CANR2X1 U11963 ( .A(mem_data1[505]), .B(n3898), .C(N8785), .D(n3659), .Z(
        n587) );
  CND3XL U11964 ( .A(n590), .B(n591), .C(n592), .Z(N9828) );
  CANR2X1 U11965 ( .A(N2580), .B(n3578), .C(n3606), .D(N7775), .Z(n592) );
  CND2X1 U11966 ( .A(N5662), .B(n3686), .Z(n591) );
  CANR2X1 U11967 ( .A(mem_data1[504]), .B(n3898), .C(N8784), .D(n3659), .Z(
        n590) );
  CND3XL U11968 ( .A(n593), .B(n594), .C(n595), .Z(N9827) );
  CANR2X1 U11969 ( .A(N2579), .B(n3578), .C(n3606), .D(N7776), .Z(n595) );
  CND2X1 U11970 ( .A(N5661), .B(n3686), .Z(n594) );
  CANR2X1 U11971 ( .A(mem_data1[503]), .B(n3898), .C(N8783), .D(n3659), .Z(
        n593) );
  CND3XL U11972 ( .A(n596), .B(n597), .C(n598), .Z(N9826) );
  CANR2X1 U11973 ( .A(N2578), .B(n3570), .C(n3606), .D(N7777), .Z(n598) );
  CND2X1 U11974 ( .A(N5660), .B(n3686), .Z(n597) );
  CANR2X1 U11975 ( .A(mem_data1[502]), .B(n3898), .C(N8782), .D(n3658), .Z(
        n596) );
  CND3XL U11976 ( .A(n599), .B(n600), .C(n601), .Z(N9825) );
  CANR2X1 U11977 ( .A(N2577), .B(n3570), .C(n3606), .D(N7778), .Z(n601) );
  CND2X1 U11978 ( .A(N5659), .B(n3686), .Z(n600) );
  CANR2X1 U11979 ( .A(mem_data1[501]), .B(n3898), .C(N8781), .D(n3658), .Z(
        n599) );
  CND3XL U11980 ( .A(n602), .B(n603), .C(n604), .Z(N9824) );
  CANR2X1 U11981 ( .A(N2576), .B(n3570), .C(n3606), .D(N7779), .Z(n604) );
  CND2X1 U11982 ( .A(N5658), .B(n3686), .Z(n603) );
  CANR2X1 U11983 ( .A(mem_data1[500]), .B(n3898), .C(N8780), .D(n3658), .Z(
        n602) );
  CND3XL U11984 ( .A(n605), .B(n606), .C(n607), .Z(N9823) );
  CND2X1 U11985 ( .A(N5657), .B(n3686), .Z(n606) );
  CANR2X1 U11986 ( .A(mem_data1[499]), .B(n3898), .C(N8779), .D(n3658), .Z(
        n605) );
  CND3XL U11987 ( .A(n608), .B(n609), .C(n610), .Z(N9822) );
  CANR2X1 U11988 ( .A(N2574), .B(n3570), .C(n3606), .D(N7781), .Z(n610) );
  CND2X1 U11989 ( .A(N5656), .B(n3686), .Z(n609) );
  CANR2X1 U11990 ( .A(mem_data1[498]), .B(n3898), .C(N8778), .D(n3658), .Z(
        n608) );
  CND3XL U11991 ( .A(n611), .B(n612), .C(n613), .Z(N9821) );
  CANR2X1 U11992 ( .A(N2573), .B(n3570), .C(n3606), .D(N7782), .Z(n613) );
  CND2X1 U11993 ( .A(N5655), .B(n3686), .Z(n612) );
  CANR2X1 U11994 ( .A(mem_data1[497]), .B(n3898), .C(N8777), .D(n3659), .Z(
        n611) );
  CND3XL U11995 ( .A(n614), .B(n615), .C(n616), .Z(N9820) );
  CND2X1 U11996 ( .A(N5654), .B(n3686), .Z(n615) );
  CANR2X1 U11997 ( .A(mem_data1[496]), .B(n3898), .C(N8776), .D(n3659), .Z(
        n614) );
  CND3XL U11998 ( .A(n617), .B(n618), .C(n619), .Z(N9819) );
  CND2X1 U11999 ( .A(N5653), .B(n3686), .Z(n618) );
  CANR2X1 U12000 ( .A(mem_data1[495]), .B(n3898), .C(N8775), .D(n3658), .Z(
        n617) );
  CND3XL U12001 ( .A(n620), .B(n621), .C(n622), .Z(N9818) );
  CND2X1 U12002 ( .A(N5652), .B(n3686), .Z(n621) );
  CANR2X1 U12003 ( .A(mem_data1[494]), .B(n3898), .C(n3644), .D(N8774), .Z(
        n620) );
  CND3XL U12004 ( .A(n641), .B(n642), .C(n643), .Z(N9811) );
  CND2X1 U12005 ( .A(N5645), .B(n3694), .Z(n642) );
  CANR2X1 U12006 ( .A(mem_data1[487]), .B(n3898), .C(n3643), .D(N8767), .Z(
        n641) );
  CND3XL U12007 ( .A(n656), .B(n657), .C(n658), .Z(N9806) );
  CND3XL U12008 ( .A(n665), .B(n666), .C(n667), .Z(N9803) );
  CND3XL U12009 ( .A(n668), .B(n669), .C(n670), .Z(N9802) );
  CND3XL U12010 ( .A(n674), .B(n675), .C(n676), .Z(N9800) );
  CND3XL U12011 ( .A(n680), .B(n681), .C(n682), .Z(N9798) );
  CND3XL U12012 ( .A(n683), .B(n684), .C(n685), .Z(N9797) );
  CND3XL U12013 ( .A(n686), .B(n687), .C(n688), .Z(N9796) );
  CND3XL U12014 ( .A(n689), .B(n690), .C(n691), .Z(N9795) );
  CND3XL U12015 ( .A(n692), .B(n693), .C(n694), .Z(N9794) );
  CND3XL U12016 ( .A(n695), .B(n696), .C(n697), .Z(N9793) );
  CND3XL U12017 ( .A(n698), .B(n699), .C(n700), .Z(N9792) );
  CND3XL U12018 ( .A(n701), .B(n702), .C(n703), .Z(N9791) );
  CND3XL U12019 ( .A(n704), .B(n705), .C(n706), .Z(N9790) );
  CND3XL U12020 ( .A(n716), .B(n717), .C(n718), .Z(N9786) );
  CND3XL U12021 ( .A(n725), .B(n726), .C(n727), .Z(N9783) );
  CND3XL U12022 ( .A(n728), .B(n729), .C(n730), .Z(N9782) );
  CND3XL U12023 ( .A(n734), .B(n735), .C(n736), .Z(N9780) );
  CND3XL U12024 ( .A(n740), .B(n741), .C(n742), .Z(N9778) );
  CND3XL U12025 ( .A(n746), .B(n747), .C(n748), .Z(N9776) );
  CND3XL U12026 ( .A(n755), .B(n756), .C(n757), .Z(N9773) );
  CANR2X1 U12027 ( .A(N2525), .B(n3571), .C(n3607), .D(N7830), .Z(n757) );
  CND2X1 U12028 ( .A(N5607), .B(n3687), .Z(n756) );
  CANR2X1 U12029 ( .A(mem_data1[449]), .B(n3898), .C(n3642), .D(N8729), .Z(
        n755) );
  CND3XL U12030 ( .A(n758), .B(n759), .C(n760), .Z(N9772) );
  CND3XL U12031 ( .A(n785), .B(n786), .C(n787), .Z(N9763) );
  CND2X1 U12032 ( .A(N5597), .B(n3687), .Z(n786) );
  CND3XL U12033 ( .A(n830), .B(n831), .C(n832), .Z(N9748) );
  CND3XL U12034 ( .A(n836), .B(n837), .C(n838), .Z(N9746) );
  CND3XL U12035 ( .A(n842), .B(n843), .C(n844), .Z(N9744) );
  CND3XL U12036 ( .A(n857), .B(n858), .C(n859), .Z(N9739) );
  CND2X1 U12037 ( .A(N5573), .B(n3689), .Z(n858) );
  CND3XL U12038 ( .A(n860), .B(n861), .C(n862), .Z(N9738) );
  CND3XL U12039 ( .A(n875), .B(n876), .C(n877), .Z(N9733) );
  CND3XL U12040 ( .A(n878), .B(n879), .C(n880), .Z(N9732) );
  CND3XL U12041 ( .A(n881), .B(n882), .C(n883), .Z(N9731) );
  CND3XL U12042 ( .A(n884), .B(n885), .C(n886), .Z(N9730) );
  CND3XL U12043 ( .A(n890), .B(n891), .C(n892), .Z(N9728) );
  CND3XL U12044 ( .A(n893), .B(n894), .C(n895), .Z(N9727) );
  CND3XL U12045 ( .A(n902), .B(n903), .C(n904), .Z(N9724) );
  CND2X1 U12046 ( .A(N5558), .B(n3684), .Z(n903) );
  CANR2X1 U12047 ( .A(mem_data1[400]), .B(n3898), .C(N8680), .D(n3659), .Z(
        n902) );
  CND3XL U12048 ( .A(n920), .B(n921), .C(n922), .Z(N9718) );
  CANR2X1 U12049 ( .A(N2470), .B(n3581), .C(n3616), .D(N7885), .Z(n922) );
  CND2X1 U12050 ( .A(N5552), .B(n3687), .Z(n921) );
  CANR2X1 U12051 ( .A(mem_data1[394]), .B(n3898), .C(N8674), .D(n3659), .Z(
        n920) );
  CND3XL U12052 ( .A(n926), .B(n927), .C(n928), .Z(N9716) );
  CND3XL U12053 ( .A(n932), .B(n933), .C(n934), .Z(N9714) );
  CND3XL U12054 ( .A(n947), .B(n948), .C(n949), .Z(N9709) );
  CND3XL U12055 ( .A(n950), .B(n951), .C(n952), .Z(N9708) );
  CANR2X1 U12056 ( .A(N2460), .B(n3582), .C(n3616), .D(N7895), .Z(n952) );
  CND3XL U12057 ( .A(n953), .B(n954), .C(n955), .Z(N9707) );
  CND3XL U12058 ( .A(n956), .B(n957), .C(n958), .Z(N9706) );
  CND3XL U12059 ( .A(n971), .B(n972), .C(n973), .Z(N9701) );
  CND2X1 U12060 ( .A(N5535), .B(n3689), .Z(n972) );
  CND3XL U12061 ( .A(n977), .B(n978), .C(n979), .Z(N9699) );
  CND2X1 U12062 ( .A(N5533), .B(n3697), .Z(n978) );
  CANR2X1 U12063 ( .A(mem_data1[375]), .B(n3898), .C(n3641), .D(N8655), .Z(
        n977) );
  CND3XL U12064 ( .A(n983), .B(n984), .C(n985), .Z(N9697) );
  CND2X1 U12065 ( .A(N5531), .B(n3689), .Z(n984) );
  CND3XL U12066 ( .A(n986), .B(n987), .C(n988), .Z(N9696) );
  CND3XL U12067 ( .A(n989), .B(n990), .C(n991), .Z(N9695) );
  CND3XL U12068 ( .A(n998), .B(n999), .C(n1000), .Z(N9692) );
  CANR2X1 U12069 ( .A(N2444), .B(n3581), .C(n3616), .D(N7911), .Z(n1000) );
  CND3XL U12070 ( .A(n1010), .B(n1011), .C(n1012), .Z(N9688) );
  CND2X1 U12071 ( .A(N5522), .B(n3698), .Z(n1011) );
  CANR2X1 U12072 ( .A(mem_data1[364]), .B(n3898), .C(N8644), .D(n3659), .Z(
        n1010) );
  CND3XL U12073 ( .A(n1022), .B(n1023), .C(n1024), .Z(N9684) );
  CND2X1 U12074 ( .A(N5518), .B(n3684), .Z(n1023) );
  CANR2X1 U12075 ( .A(mem_data1[360]), .B(n3898), .C(N8640), .D(n3659), .Z(
        n1022) );
  CND3XL U12076 ( .A(n1088), .B(n1089), .C(n1090), .Z(N9662) );
  CND3XL U12077 ( .A(n1094), .B(n1095), .C(n1096), .Z(N9660) );
  CND3XL U12078 ( .A(n1100), .B(n1101), .C(n1102), .Z(N9658) );
  CND3XL U12079 ( .A(n1103), .B(n1104), .C(n1105), .Z(N9657) );
  CND3XL U12080 ( .A(n1106), .B(n1107), .C(n1108), .Z(N9656) );
  CND3XL U12081 ( .A(n1109), .B(n1110), .C(n1111), .Z(N9655) );
  CND3XL U12082 ( .A(n1112), .B(n1113), .C(n1114), .Z(N9654) );
  CND3XL U12083 ( .A(n1115), .B(n1116), .C(n1117), .Z(N9653) );
  CND3XL U12084 ( .A(n1118), .B(n1119), .C(n1120), .Z(N9652) );
  CND3XL U12085 ( .A(n1136), .B(n1137), .C(n1138), .Z(N9646) );
  CND3XL U12086 ( .A(n1145), .B(n1146), .C(n1147), .Z(N9643) );
  CND3XL U12087 ( .A(n1148), .B(n1149), .C(n1150), .Z(N9642) );
  CND3XL U12088 ( .A(n1166), .B(n1167), .C(n1168), .Z(N9636) );
  CND3XL U12089 ( .A(n1169), .B(n1170), .C(n1171), .Z(N9635) );
  CND3XL U12090 ( .A(n1172), .B(n1173), .C(n1174), .Z(N9634) );
  CND3XL U12091 ( .A(n1178), .B(n1179), .C(n1180), .Z(N9632) );
  CND3XL U12092 ( .A(n1181), .B(n1182), .C(n1183), .Z(N9631) );
  CND3XL U12093 ( .A(n1184), .B(n1185), .C(n1186), .Z(N9630) );
  CND2X1 U12094 ( .A(N5464), .B(n3696), .Z(n1185) );
  CANR2X1 U12095 ( .A(mem_data1[306]), .B(n3898), .C(n3640), .D(N8586), .Z(
        n1184) );
  CND3XL U12096 ( .A(n1196), .B(n1197), .C(n1198), .Z(N9626) );
  CND2X1 U12097 ( .A(N5460), .B(n3693), .Z(n1197) );
  CANR2X1 U12098 ( .A(mem_data1[302]), .B(n3898), .C(n3640), .D(N8582), .Z(
        n1196) );
  CND3XL U12099 ( .A(n1205), .B(n1206), .C(n1207), .Z(N9623) );
  CND2X1 U12100 ( .A(N5457), .B(n3690), .Z(n1206) );
  CND3XL U12101 ( .A(n1235), .B(n1236), .C(n1237), .Z(N9613) );
  CND3XL U12102 ( .A(n1238), .B(n1239), .C(n1240), .Z(N9612) );
  CANR2X1 U12103 ( .A(N2364), .B(n3582), .C(n3617), .D(N7991), .Z(n1240) );
  CND2X1 U12104 ( .A(N5446), .B(n3696), .Z(n1239) );
  CANR2X1 U12105 ( .A(mem_data1[288]), .B(n3898), .C(n3640), .D(N8568), .Z(
        n1238) );
  CND3XL U12106 ( .A(n1241), .B(n1242), .C(n1243), .Z(N9611) );
  CND2X1 U12107 ( .A(N5445), .B(n3696), .Z(n1242) );
  CANR2X1 U12108 ( .A(mem_data1[287]), .B(n3898), .C(n3640), .D(N8567), .Z(
        n1241) );
  CND3XL U12109 ( .A(n1247), .B(n1248), .C(n1249), .Z(N9609) );
  CND2X1 U12110 ( .A(N5443), .B(n3684), .Z(n1248) );
  CANR2X1 U12111 ( .A(mem_data1[285]), .B(n3898), .C(n3640), .D(N8565), .Z(
        n1247) );
  CND3XL U12112 ( .A(n1250), .B(n1251), .C(n1252), .Z(N9608) );
  CANR2X1 U12113 ( .A(N2360), .B(n3585), .C(n3622), .D(N7995), .Z(n1252) );
  CND2X1 U12114 ( .A(N5442), .B(n3697), .Z(n1251) );
  CANR2X1 U12115 ( .A(mem_data1[284]), .B(n3898), .C(n3640), .D(N8564), .Z(
        n1250) );
  CND3XL U12116 ( .A(n1256), .B(n1257), .C(n1258), .Z(N9606) );
  CND3XL U12117 ( .A(n1259), .B(n1260), .C(n1261), .Z(N9605) );
  CANR2X1 U12118 ( .A(N2357), .B(n3585), .C(n3620), .D(N7998), .Z(n1261) );
  CND2X1 U12119 ( .A(N5439), .B(n3685), .Z(n1260) );
  CANR2X1 U12120 ( .A(mem_data1[281]), .B(n3898), .C(n3640), .D(N8561), .Z(
        n1259) );
  CND3XL U12121 ( .A(n1262), .B(n1263), .C(n1264), .Z(N9604) );
  CANR2X1 U12122 ( .A(N2356), .B(n3585), .C(n3620), .D(N7999), .Z(n1264) );
  CND2X1 U12123 ( .A(N5438), .B(n3683), .Z(n1263) );
  CANR2X1 U12124 ( .A(mem_data1[280]), .B(n3898), .C(n3640), .D(N8560), .Z(
        n1262) );
  CND3XL U12125 ( .A(n1274), .B(n1275), .C(n1276), .Z(N9600) );
  CANR2X1 U12126 ( .A(N2352), .B(n3586), .C(n3620), .D(N8003), .Z(n1276) );
  CND2X1 U12127 ( .A(N5434), .B(n3686), .Z(n1275) );
  CANR2X1 U12128 ( .A(mem_data1[276]), .B(n3898), .C(n3640), .D(N8556), .Z(
        n1274) );
  CND3XL U12129 ( .A(n1277), .B(n1278), .C(n1279), .Z(N9599) );
  CND2X1 U12130 ( .A(N5433), .B(n3685), .Z(n1278) );
  CANR2X1 U12131 ( .A(mem_data1[275]), .B(n3898), .C(n3640), .D(N8555), .Z(
        n1277) );
  CND3XL U12132 ( .A(n1280), .B(n1281), .C(n1282), .Z(N9598) );
  CANR2X1 U12133 ( .A(N2350), .B(n3586), .C(n3620), .D(N8005), .Z(n1282) );
  CND2X1 U12134 ( .A(N5432), .B(n3688), .Z(n1281) );
  CANR2X1 U12135 ( .A(mem_data1[274]), .B(n3898), .C(n3640), .D(N8554), .Z(
        n1280) );
  CND3XL U12136 ( .A(n1286), .B(n1287), .C(n1288), .Z(N9596) );
  CANR2X1 U12137 ( .A(N2348), .B(n3586), .C(n3620), .D(N8007), .Z(n1288) );
  CND2X1 U12138 ( .A(N5430), .B(n3689), .Z(n1287) );
  CANR2X1 U12139 ( .A(mem_data1[272]), .B(n3898), .C(n3640), .D(N8552), .Z(
        n1286) );
  CND3XL U12140 ( .A(n1292), .B(n1293), .C(n1294), .Z(N9594) );
  CANR2X1 U12141 ( .A(N2346), .B(n3586), .C(n3621), .D(N8009), .Z(n1294) );
  CND2X1 U12142 ( .A(N5428), .B(n3695), .Z(n1293) );
  CANR2X1 U12143 ( .A(mem_data1[270]), .B(n3898), .C(n3640), .D(N8550), .Z(
        n1292) );
  CND3XL U12144 ( .A(n1295), .B(n1296), .C(n1297), .Z(N9593) );
  CND2X1 U12145 ( .A(N5427), .B(n3691), .Z(n1296) );
  CANR2X1 U12146 ( .A(mem_data1[269]), .B(n3898), .C(n3640), .D(N8549), .Z(
        n1295) );
  CND3XL U12147 ( .A(n1298), .B(n1299), .C(n1300), .Z(N9592) );
  CANR2X1 U12148 ( .A(N2344), .B(n3586), .C(n3621), .D(N8011), .Z(n1300) );
  CND2X1 U12149 ( .A(N5426), .B(n3693), .Z(n1299) );
  CANR2X1 U12150 ( .A(mem_data1[268]), .B(n3898), .C(n3640), .D(N8548), .Z(
        n1298) );
  CND3XL U12151 ( .A(n1301), .B(n1302), .C(n1303), .Z(N9591) );
  CND2X1 U12152 ( .A(N5425), .B(n3683), .Z(n1302) );
  CANR2X1 U12153 ( .A(mem_data1[267]), .B(n3898), .C(n3640), .D(N8547), .Z(
        n1301) );
  CND3XL U12154 ( .A(n1304), .B(n1305), .C(n1306), .Z(N9590) );
  CANR2X1 U12155 ( .A(N2342), .B(n3586), .C(n3621), .D(N8013), .Z(n1306) );
  CND2X1 U12156 ( .A(N5424), .B(n3684), .Z(n1305) );
  CANR2X1 U12157 ( .A(mem_data1[266]), .B(n3898), .C(n3640), .D(N8546), .Z(
        n1304) );
  CND3XL U12158 ( .A(n1307), .B(n1308), .C(n1309), .Z(N9589) );
  CANR2X1 U12159 ( .A(N2341), .B(n3586), .C(n3621), .D(N8014), .Z(n1309) );
  CND2X1 U12160 ( .A(N5423), .B(n3696), .Z(n1308) );
  CANR2X1 U12161 ( .A(mem_data1[265]), .B(n3898), .C(n3640), .D(N8545), .Z(
        n1307) );
  CND3XL U12162 ( .A(n1310), .B(n1311), .C(n1312), .Z(N9588) );
  CND3XL U12163 ( .A(n1313), .B(n1314), .C(n1315), .Z(N9587) );
  CND3XL U12164 ( .A(n1316), .B(n1317), .C(n1318), .Z(N9586) );
  CANR2X1 U12165 ( .A(N2338), .B(n3586), .C(n3621), .D(N8017), .Z(n1318) );
  CND2X1 U12166 ( .A(N5420), .B(n3694), .Z(n1317) );
  CANR2X1 U12167 ( .A(mem_data1[262]), .B(n3898), .C(n3640), .D(N8542), .Z(
        n1316) );
  CND3XL U12168 ( .A(n1322), .B(n1323), .C(n1324), .Z(N9584) );
  CND3XL U12169 ( .A(n1328), .B(n1329), .C(n1330), .Z(N9582) );
  CND3XL U12170 ( .A(n1337), .B(n1338), .C(n1339), .Z(N9579) );
  CND3XL U12171 ( .A(n1340), .B(n1341), .C(n1342), .Z(N9578) );
  CND3XL U12172 ( .A(n1361), .B(n1362), .C(n1363), .Z(N9571) );
  CND2X1 U12173 ( .A(N5405), .B(n3683), .Z(n1362) );
  CANR2X1 U12174 ( .A(mem_data1[247]), .B(n3898), .C(N8527), .D(n3659), .Z(
        n1361) );
  CND3XL U12175 ( .A(n1370), .B(n1371), .C(n1372), .Z(N9568) );
  CND2X1 U12176 ( .A(N5402), .B(n3687), .Z(n1371) );
  CANR2X1 U12177 ( .A(mem_data1[244]), .B(n3898), .C(N8524), .D(n3659), .Z(
        n1370) );
  CND3XL U12178 ( .A(n1379), .B(n1380), .C(n1381), .Z(N9565) );
  CND3XL U12179 ( .A(n1382), .B(n1383), .C(n1384), .Z(N9564) );
  CND3XL U12180 ( .A(n1385), .B(n1386), .C(n1387), .Z(N9563) );
  CND3XL U12181 ( .A(n1388), .B(n1389), .C(n1390), .Z(N9562) );
  CND2X1 U12182 ( .A(N5396), .B(n3695), .Z(n1389) );
  CND3XL U12183 ( .A(n1391), .B(n1392), .C(n1393), .Z(N9561) );
  CND3XL U12184 ( .A(n1394), .B(n1395), .C(n1396), .Z(N9560) );
  CND3XL U12185 ( .A(n1397), .B(n1398), .C(n1399), .Z(N9559) );
  CND3XL U12186 ( .A(n1400), .B(n1401), .C(n1402), .Z(N9558) );
  CND3XL U12187 ( .A(n1403), .B(n1404), .C(n1405), .Z(N9557) );
  CND3XL U12188 ( .A(n1406), .B(n1407), .C(n1408), .Z(N9556) );
  CND3XL U12189 ( .A(n1409), .B(n1410), .C(n1411), .Z(N9555) );
  CND3XL U12190 ( .A(n1412), .B(n1413), .C(n1414), .Z(N9554) );
  CND2X1 U12191 ( .A(N5388), .B(n3698), .Z(n1413) );
  CND3XL U12192 ( .A(n1415), .B(n1416), .C(n1417), .Z(N9553) );
  CND3XL U12193 ( .A(n1418), .B(n1419), .C(n1420), .Z(N9552) );
  CND3XL U12194 ( .A(n1421), .B(n1422), .C(n1423), .Z(N9551) );
  CND3XL U12195 ( .A(n1424), .B(n1425), .C(n1426), .Z(N9550) );
  CND3XL U12196 ( .A(n1427), .B(n1428), .C(n1429), .Z(N9549) );
  CND3XL U12197 ( .A(n1430), .B(n1431), .C(n1432), .Z(N9548) );
  CND3XL U12198 ( .A(n1433), .B(n1434), .C(n1435), .Z(N9547) );
  CND3XL U12199 ( .A(n1436), .B(n1437), .C(n1438), .Z(N9546) );
  CND2X1 U12200 ( .A(N5380), .B(n3698), .Z(n1437) );
  CANR2X1 U12201 ( .A(mem_data1[222]), .B(n3898), .C(N8502), .D(n3647), .Z(
        n1436) );
  CND3XL U12202 ( .A(n1439), .B(n1440), .C(n1441), .Z(N9545) );
  CANR2X1 U12203 ( .A(N2297), .B(n3579), .C(n3621), .D(N8058), .Z(n1441) );
  CND2X1 U12204 ( .A(N5379), .B(n3697), .Z(n1440) );
  CANR2X1 U12205 ( .A(mem_data1[221]), .B(n3898), .C(N8501), .D(n3649), .Z(
        n1439) );
  CND3XL U12206 ( .A(n1445), .B(n1446), .C(n1447), .Z(N9543) );
  CND3XL U12207 ( .A(n1448), .B(n1449), .C(n1450), .Z(N9542) );
  CND3XL U12208 ( .A(n1451), .B(n1452), .C(n1453), .Z(N9541) );
  CND3XL U12209 ( .A(n1454), .B(n1455), .C(n1456), .Z(N9540) );
  CND3XL U12210 ( .A(n1457), .B(n1458), .C(n1459), .Z(N9539) );
  CND3XL U12211 ( .A(n1460), .B(n1461), .C(n1462), .Z(N9538) );
  CND3XL U12212 ( .A(n1463), .B(n1464), .C(n1465), .Z(N9537) );
  CND3XL U12213 ( .A(n1466), .B(n1467), .C(n1468), .Z(N9536) );
  CND3XL U12214 ( .A(n1469), .B(n1470), .C(n1471), .Z(N9535) );
  CND3XL U12215 ( .A(n1472), .B(n1473), .C(n1474), .Z(N9534) );
  CND3XL U12216 ( .A(n1475), .B(n1476), .C(n1477), .Z(N9533) );
  CND3XL U12217 ( .A(n1478), .B(n1479), .C(n1480), .Z(N9532) );
  CND3XL U12218 ( .A(n1481), .B(n1482), .C(n1483), .Z(N9531) );
  CND3XL U12219 ( .A(n1484), .B(n1485), .C(n1486), .Z(N9530) );
  CND3XL U12220 ( .A(n1487), .B(n1488), .C(n1489), .Z(N9529) );
  CND3XL U12221 ( .A(n1490), .B(n1491), .C(n1492), .Z(N9528) );
  CND3XL U12222 ( .A(n1493), .B(n1494), .C(n1495), .Z(N9527) );
  CND3XL U12223 ( .A(n1496), .B(n1497), .C(n1498), .Z(N9526) );
  CND3XL U12224 ( .A(n1499), .B(n1500), .C(n1501), .Z(N9525) );
  CND3XL U12225 ( .A(n1502), .B(n1503), .C(n1504), .Z(N9524) );
  CND3XL U12226 ( .A(n1505), .B(n1506), .C(n1507), .Z(N9523) );
  CANR2X1 U12227 ( .A(N2275), .B(n3580), .C(n3614), .D(N8080), .Z(n1507) );
  CND2X1 U12228 ( .A(N5357), .B(n3694), .Z(n1506) );
  CANR2X1 U12229 ( .A(mem_data1[199]), .B(n3898), .C(N8479), .D(n3650), .Z(
        n1505) );
  CND3XL U12230 ( .A(n1508), .B(n1509), .C(n1510), .Z(N9522) );
  CND3XL U12231 ( .A(n1511), .B(n1512), .C(n1513), .Z(N9521) );
  CND3XL U12232 ( .A(n1514), .B(n1515), .C(n1516), .Z(N9520) );
  CND3XL U12233 ( .A(n1517), .B(n1518), .C(n1519), .Z(N9519) );
  CND3XL U12234 ( .A(n1520), .B(n1521), .C(n1522), .Z(N9518) );
  CND3XL U12235 ( .A(n1523), .B(n1524), .C(n1525), .Z(N9517) );
  CND3XL U12236 ( .A(n1526), .B(n1527), .C(n1528), .Z(N9516) );
  CND3XL U12237 ( .A(n1529), .B(n1530), .C(n1531), .Z(N9515) );
  CND3XL U12238 ( .A(n1532), .B(n1533), .C(n1534), .Z(N9514) );
  CND3XL U12239 ( .A(n1538), .B(n1539), .C(n1540), .Z(N9512) );
  CND3XL U12240 ( .A(n1550), .B(n1551), .C(n1552), .Z(N9508) );
  CND3XL U12241 ( .A(n1562), .B(n1563), .C(n1564), .Z(N9504) );
  CND3XL U12242 ( .A(n1565), .B(n1566), .C(n1567), .Z(N9503) );
  CND3XL U12243 ( .A(n1568), .B(n1569), .C(n1570), .Z(N9502) );
  CND3XL U12244 ( .A(n1571), .B(n1572), .C(n1573), .Z(N9501) );
  CND3XL U12245 ( .A(n1574), .B(n1575), .C(n1576), .Z(N9500) );
  CND3XL U12246 ( .A(n1577), .B(n1578), .C(n1579), .Z(N9499) );
  CND3XL U12247 ( .A(n1580), .B(n1581), .C(n1582), .Z(N9498) );
  CND3XL U12248 ( .A(n1583), .B(n1584), .C(n1585), .Z(N9497) );
  CND3XL U12249 ( .A(n1586), .B(n1587), .C(n1588), .Z(N9496) );
  CND3XL U12250 ( .A(n1589), .B(n1590), .C(n1591), .Z(N9495) );
  CND3XL U12251 ( .A(n1592), .B(n1593), .C(n1594), .Z(N9494) );
  CND3XL U12252 ( .A(n1595), .B(n1596), .C(n1597), .Z(N9493) );
  CND3XL U12253 ( .A(n1598), .B(n1599), .C(n1600), .Z(N9492) );
  CND3XL U12254 ( .A(n1601), .B(n1602), .C(n1603), .Z(N9491) );
  CND3XL U12255 ( .A(n1604), .B(n1605), .C(n1606), .Z(N9490) );
  CND3XL U12256 ( .A(n1607), .B(n1608), .C(n1609), .Z(N9489) );
  CND3XL U12257 ( .A(n1610), .B(n1611), .C(n1612), .Z(N9488) );
  CND3XL U12258 ( .A(n1613), .B(n1614), .C(n1615), .Z(N9487) );
  CND3XL U12259 ( .A(n1616), .B(n1617), .C(n1618), .Z(N9486) );
  CND2X1 U12260 ( .A(N5320), .B(n3695), .Z(n1617) );
  CND3XL U12261 ( .A(n1619), .B(n1620), .C(n1621), .Z(N9485) );
  CND3XL U12262 ( .A(n1622), .B(n1623), .C(n1624), .Z(N9484) );
  CND3XL U12263 ( .A(n1625), .B(n1626), .C(n1627), .Z(N9483) );
  CND3XL U12264 ( .A(n1628), .B(n1629), .C(n1630), .Z(N9482) );
  CND3XL U12265 ( .A(n1631), .B(n1632), .C(n1633), .Z(N9481) );
  CND3XL U12266 ( .A(n1634), .B(n1635), .C(n1636), .Z(N9480) );
  CND3XL U12267 ( .A(n1637), .B(n1638), .C(n1639), .Z(N9479) );
  CND3XL U12268 ( .A(n1640), .B(n1641), .C(n1642), .Z(N9478) );
  CND3XL U12269 ( .A(n1643), .B(n1644), .C(n1645), .Z(N9477) );
  CND3XL U12270 ( .A(n1646), .B(n1647), .C(n1648), .Z(N9476) );
  CND3XL U12271 ( .A(n1649), .B(n1650), .C(n1651), .Z(N9475) );
  CND3XL U12272 ( .A(n1652), .B(n1653), .C(n1654), .Z(N9474) );
  CND3XL U12273 ( .A(n1655), .B(n1656), .C(n1657), .Z(N9473) );
  CND3XL U12274 ( .A(n1658), .B(n1659), .C(n1660), .Z(N9472) );
  CND3XL U12275 ( .A(n1661), .B(n1662), .C(n1663), .Z(N9471) );
  CND3XL U12276 ( .A(n1664), .B(n1665), .C(n1666), .Z(N9470) );
  CND3XL U12277 ( .A(n1667), .B(n1668), .C(n1669), .Z(N9469) );
  CND3XL U12278 ( .A(n1670), .B(n1671), .C(n1672), .Z(N9468) );
  CND3XL U12279 ( .A(n1673), .B(n1674), .C(n1675), .Z(N9467) );
  CND3XL U12280 ( .A(n1676), .B(n1677), .C(n1678), .Z(N9466) );
  CND3XL U12281 ( .A(n1679), .B(n1680), .C(n1681), .Z(N9465) );
  CND3XL U12282 ( .A(n1682), .B(n1683), .C(n1684), .Z(N9464) );
  CND3XL U12283 ( .A(n1685), .B(n1686), .C(n1687), .Z(N9463) );
  CND3XL U12284 ( .A(n1688), .B(n1689), .C(n1690), .Z(N9462) );
  CND3XL U12285 ( .A(n1691), .B(n1692), .C(n1693), .Z(N9461) );
  CND3XL U12286 ( .A(n1694), .B(n1695), .C(n1696), .Z(N9460) );
  CND3XL U12287 ( .A(n1697), .B(n1698), .C(n1699), .Z(N9459) );
  CND3XL U12288 ( .A(n1700), .B(n1701), .C(n1702), .Z(N9458) );
  CND3XL U12289 ( .A(n1703), .B(n1704), .C(n1705), .Z(N9457) );
  CND3XL U12290 ( .A(n1706), .B(n1707), .C(n1708), .Z(N9456) );
  CND3XL U12291 ( .A(n1709), .B(n1710), .C(n1711), .Z(N9455) );
  CND3XL U12292 ( .A(n1712), .B(n1713), .C(n1714), .Z(N9454) );
  CND3XL U12293 ( .A(n1715), .B(n1716), .C(n1717), .Z(N9453) );
  CND3XL U12294 ( .A(n1718), .B(n1719), .C(n1720), .Z(N9452) );
  CANR2X1 U12295 ( .A(N2204), .B(n3588), .C(n3623), .D(N8151), .Z(n1720) );
  CND3XL U12296 ( .A(n1721), .B(n1722), .C(n1723), .Z(N9451) );
  CND3XL U12297 ( .A(n1724), .B(n1725), .C(n1726), .Z(N9450) );
  CND3XL U12298 ( .A(n1727), .B(n1728), .C(n1729), .Z(N9449) );
  CND3XL U12299 ( .A(n1730), .B(n1731), .C(n1732), .Z(N9448) );
  CND3XL U12300 ( .A(n1733), .B(n1734), .C(n1735), .Z(N9447) );
  CND2X1 U12301 ( .A(N5281), .B(n3697), .Z(n1734) );
  CND3XL U12302 ( .A(n1736), .B(n1737), .C(n1738), .Z(N9446) );
  CND3XL U12303 ( .A(n1739), .B(n1740), .C(n1741), .Z(N9445) );
  CND3XL U12304 ( .A(n1745), .B(n1746), .C(n1747), .Z(N9443) );
  CND2X1 U12305 ( .A(N5277), .B(n3697), .Z(n1746) );
  CND3XL U12306 ( .A(n1751), .B(n1752), .C(n1753), .Z(N9441) );
  CANR2X1 U12307 ( .A(N2193), .B(n3589), .C(n3623), .D(N8162), .Z(n1753) );
  CND2X1 U12308 ( .A(N5275), .B(n3697), .Z(n1752) );
  CANR2X1 U12309 ( .A(mem_data1[117]), .B(n3898), .C(N8397), .D(n3646), .Z(
        n1751) );
  CND3XL U12310 ( .A(n1757), .B(n1758), .C(n1759), .Z(N9439) );
  CND2X1 U12311 ( .A(N5273), .B(n3696), .Z(n1758) );
  CND3XL U12312 ( .A(n1760), .B(n1761), .C(n1762), .Z(N9438) );
  CND3XL U12313 ( .A(n1766), .B(n1767), .C(n1768), .Z(N9436) );
  CND3XL U12314 ( .A(n1772), .B(n1773), .C(n1774), .Z(N9434) );
  CND2X1 U12315 ( .A(N5268), .B(n3697), .Z(n1773) );
  CND3XL U12316 ( .A(n1775), .B(n1776), .C(n1777), .Z(N9433) );
  CND3XL U12317 ( .A(n1778), .B(n1779), .C(n1780), .Z(N9432) );
  CND3XL U12318 ( .A(n1781), .B(n1782), .C(n1783), .Z(N9431) );
  CND3XL U12319 ( .A(n1784), .B(n1785), .C(n1786), .Z(N9430) );
  CND3XL U12320 ( .A(n1787), .B(n1788), .C(n1789), .Z(N9429) );
  CND3XL U12321 ( .A(n1790), .B(n1791), .C(n1792), .Z(N9428) );
  CND3XL U12322 ( .A(n1793), .B(n1794), .C(n1795), .Z(N9427) );
  CND3XL U12323 ( .A(n1796), .B(n1797), .C(n1798), .Z(N9426) );
  CND2X1 U12324 ( .A(N5260), .B(n3688), .Z(n1797) );
  CND3XL U12325 ( .A(n1799), .B(n1800), .C(n1801), .Z(N9425) );
  CND3XL U12326 ( .A(n1802), .B(n1803), .C(n1804), .Z(N9424) );
  CND3XL U12327 ( .A(n1805), .B(n1806), .C(n1807), .Z(N9423) );
  CND3XL U12328 ( .A(n1808), .B(n1809), .C(n1810), .Z(N9422) );
  CND3XL U12329 ( .A(n1811), .B(n1812), .C(n1813), .Z(N9421) );
  CND3XL U12330 ( .A(n1814), .B(n1815), .C(n1816), .Z(N9420) );
  CANR2X1 U12331 ( .A(N2172), .B(n3590), .C(n3623), .D(N8183), .Z(n1816) );
  CND3XL U12332 ( .A(n1817), .B(n1818), .C(n1819), .Z(N9419) );
  CND3XL U12333 ( .A(n1820), .B(n1821), .C(n1822), .Z(N9418) );
  CND2X1 U12334 ( .A(N5252), .B(n3685), .Z(n1821) );
  CND3XL U12335 ( .A(n1823), .B(n1824), .C(n1825), .Z(N9417) );
  CND3XL U12336 ( .A(n1826), .B(n1827), .C(n1828), .Z(N9416) );
  CND3XL U12337 ( .A(n1829), .B(n1830), .C(n1831), .Z(N9415) );
  CND3XL U12338 ( .A(n1832), .B(n1833), .C(n1834), .Z(N9414) );
  CND3XL U12339 ( .A(n1835), .B(n1836), .C(n1837), .Z(N9413) );
  CANR2X1 U12340 ( .A(N2165), .B(n3590), .C(n3625), .D(N8190), .Z(n1837) );
  CND2X1 U12341 ( .A(N5247), .B(n3690), .Z(n1836) );
  CANR2X1 U12342 ( .A(mem_data1[89]), .B(n3898), .C(N8369), .D(n3645), .Z(
        n1835) );
  CND3XL U12343 ( .A(n1838), .B(n1839), .C(n1840), .Z(N9412) );
  CND3XL U12344 ( .A(n1841), .B(n1842), .C(n1843), .Z(N9411) );
  CND3XL U12345 ( .A(n1844), .B(n1845), .C(n1846), .Z(N9410) );
  CND3XL U12346 ( .A(n1847), .B(n1848), .C(n1849), .Z(N9409) );
  CND3XL U12347 ( .A(n1850), .B(n1851), .C(n1852), .Z(N9408) );
  CND3XL U12348 ( .A(n1853), .B(n1854), .C(n1855), .Z(N9407) );
  CND3XL U12349 ( .A(n1856), .B(n1857), .C(n1858), .Z(N9406) );
  CND3XL U12350 ( .A(n1859), .B(n1860), .C(n1861), .Z(N9405) );
  CND3XL U12351 ( .A(n1862), .B(n1863), .C(n1864), .Z(N9404) );
  CND3XL U12352 ( .A(n1865), .B(n1866), .C(n1867), .Z(N9403) );
  CND3XL U12353 ( .A(n1868), .B(n1869), .C(n1870), .Z(N9402) );
  CND3XL U12354 ( .A(n1871), .B(n1872), .C(n1873), .Z(N9401) );
  CND3XL U12355 ( .A(n1874), .B(n1875), .C(n1876), .Z(N9400) );
  CND3XL U12356 ( .A(n1877), .B(n1878), .C(n1879), .Z(N9399) );
  CND3XL U12357 ( .A(n1880), .B(n1881), .C(n1882), .Z(N9398) );
  CND3XL U12358 ( .A(n1883), .B(n1884), .C(n1885), .Z(N9397) );
  CND3XL U12359 ( .A(n1886), .B(n1887), .C(n1888), .Z(N9396) );
  CND3XL U12360 ( .A(n1889), .B(n1890), .C(n1891), .Z(N9395) );
  CND3XL U12361 ( .A(n1892), .B(n1893), .C(n1894), .Z(N9394) );
  CND3XL U12362 ( .A(n1895), .B(n1896), .C(n1897), .Z(N9393) );
  CND3XL U12363 ( .A(n1898), .B(n1899), .C(n1900), .Z(N9392) );
  CND3XL U12364 ( .A(n1901), .B(n1902), .C(n1903), .Z(N9391) );
  CND3XL U12365 ( .A(n1904), .B(n1905), .C(n1906), .Z(N9390) );
  CND3XL U12366 ( .A(n1907), .B(n1908), .C(n1909), .Z(N9389) );
  CND3XL U12367 ( .A(n1910), .B(n1911), .C(n1912), .Z(N9388) );
  CANR2X1 U12368 ( .A(N2140), .B(n3590), .C(n3624), .D(N8215), .Z(n1912) );
  CND3XL U12369 ( .A(n1913), .B(n1914), .C(n1915), .Z(N9387) );
  CND3XL U12370 ( .A(n1916), .B(n1917), .C(n1918), .Z(N9386) );
  CND3XL U12371 ( .A(n1922), .B(n1923), .C(n1924), .Z(N9384) );
  CND3XL U12372 ( .A(n1931), .B(n1932), .C(n1933), .Z(N9381) );
  CND3XL U12373 ( .A(n1934), .B(n1935), .C(n1936), .Z(N9380) );
  CND3XL U12374 ( .A(n1937), .B(n1938), .C(n1939), .Z(N9379) );
  CND3XL U12375 ( .A(n1940), .B(n1941), .C(n1942), .Z(N9378) );
  CND3XL U12376 ( .A(n1943), .B(n1944), .C(n1945), .Z(N9377) );
  CND3XL U12377 ( .A(n1946), .B(n1947), .C(n1948), .Z(N9376) );
  CND3XL U12378 ( .A(n1949), .B(n1950), .C(n1951), .Z(N9375) );
  CND3XL U12379 ( .A(n1952), .B(n1953), .C(n1954), .Z(N9374) );
  CND3XL U12380 ( .A(n1955), .B(n1956), .C(n1957), .Z(N9373) );
  CND3XL U12381 ( .A(n1958), .B(n1959), .C(n1960), .Z(N9372) );
  CND3XL U12382 ( .A(n1961), .B(n1962), .C(n1963), .Z(N9371) );
  CND3XL U12383 ( .A(n1964), .B(n1965), .C(n1966), .Z(N9370) );
  CND3XL U12384 ( .A(n1967), .B(n1968), .C(n1969), .Z(N9369) );
  CND3XL U12385 ( .A(n1970), .B(n1971), .C(n1972), .Z(N9368) );
  CND3XL U12386 ( .A(n1973), .B(n1974), .C(n1975), .Z(N9367) );
  CND3XL U12387 ( .A(n1976), .B(n1977), .C(n1978), .Z(N9366) );
  CND3XL U12388 ( .A(n1979), .B(n1980), .C(n1981), .Z(N9365) );
  CND3XL U12389 ( .A(n1982), .B(n1983), .C(n1984), .Z(N9364) );
  CND3XL U12390 ( .A(n1985), .B(n1986), .C(n1987), .Z(N9363) );
  CND3XL U12391 ( .A(n1988), .B(n1989), .C(n1990), .Z(N9362) );
  CND3XL U12392 ( .A(n1991), .B(n1992), .C(n1993), .Z(N9361) );
  CND3XL U12393 ( .A(n1994), .B(n1995), .C(n1996), .Z(N9360) );
  CND3XL U12394 ( .A(n1997), .B(n1998), .C(n1999), .Z(N9359) );
  CND3XL U12395 ( .A(n2000), .B(n2001), .C(n2002), .Z(N9358) );
  CND3XL U12396 ( .A(n2003), .B(n2004), .C(n2005), .Z(N9357) );
  CND3XL U12397 ( .A(n2006), .B(n2007), .C(n2008), .Z(N9356) );
  CND3XL U12398 ( .A(n2009), .B(n2010), .C(n2011), .Z(N9355) );
  CND3XL U12399 ( .A(n2012), .B(n2013), .C(n2014), .Z(N9354) );
  CND3XL U12400 ( .A(n2015), .B(n2016), .C(n2017), .Z(N9353) );
  CND3XL U12401 ( .A(n2018), .B(n2019), .C(n2020), .Z(N9352) );
  CND3XL U12402 ( .A(n2021), .B(n2022), .C(n2023), .Z(N9351) );
  CND3XL U12403 ( .A(n2024), .B(n2025), .C(n2026), .Z(N9350) );
  CND3XL U12404 ( .A(n2027), .B(n2028), .C(n2029), .Z(N9349) );
  CND3XL U12405 ( .A(n2030), .B(n2031), .C(n2032), .Z(N9348) );
  CND3XL U12406 ( .A(n2033), .B(n2034), .C(n2035), .Z(N9347) );
  CND3XL U12407 ( .A(n2036), .B(n2037), .C(n2038), .Z(N9346) );
  CND3XL U12408 ( .A(n2039), .B(n2040), .C(n2041), .Z(N9345) );
  CND3XL U12409 ( .A(n2042), .B(n2043), .C(n2044), .Z(N9344) );
  CND3XL U12410 ( .A(n2045), .B(n2046), .C(n2047), .Z(N9343) );
  CND3XL U12411 ( .A(n2048), .B(n2049), .C(n2050), .Z(N9342) );
  CND3XL U12412 ( .A(n2051), .B(n2052), .C(n2053), .Z(N9341) );
  CND3XL U12413 ( .A(n2054), .B(n2055), .C(n2056), .Z(N9340) );
  CND3XL U12414 ( .A(n2057), .B(n2058), .C(n2059), .Z(N9339) );
  CND3XL U12415 ( .A(n2060), .B(n2061), .C(n2062), .Z(N9338) );
  CND3XL U12416 ( .A(n2063), .B(n2064), .C(n2065), .Z(N9337) );
  CND3XL U12417 ( .A(n2066), .B(n2067), .C(n2068), .Z(N9336) );
  CND3XL U12418 ( .A(n2069), .B(n2070), .C(n2071), .Z(N9335) );
  CND3XL U12419 ( .A(n2072), .B(n2073), .C(n2074), .Z(N9334) );
  CND3XL U12420 ( .A(n2075), .B(n2076), .C(n2077), .Z(N9333) );
  CND3XL U12421 ( .A(n2078), .B(n2079), .C(n2080), .Z(N9332) );
  CND3XL U12422 ( .A(n2081), .B(n2082), .C(n2083), .Z(N9331) );
  CND3XL U12423 ( .A(n2084), .B(n2085), .C(n2086), .Z(N9330) );
  CANR2X1 U12424 ( .A(N2082), .B(n3593), .C(n3626), .D(N8273), .Z(n2086) );
  CND3XL U12425 ( .A(n2087), .B(n2088), .C(n2089), .Z(N9329) );
  CANR2X1 U12426 ( .A(N2081), .B(n3593), .C(n3626), .D(N8274), .Z(n2089) );
  CND3XL U12427 ( .A(n2093), .B(n2094), .C(n2095), .Z(N9327) );
  CANR2X1 U12428 ( .A(N2079), .B(n3593), .C(n3628), .D(N8276), .Z(n2095) );
  CND3XL U12429 ( .A(n2096), .B(n2097), .C(n2098), .Z(N9326) );
  CANR2X1 U12430 ( .A(N2078), .B(n3592), .C(n3626), .D(N8277), .Z(n2098) );
  CND3XL U12431 ( .A(n2099), .B(n2100), .C(n2101), .Z(N9325) );
  CANR2X1 U12432 ( .A(N2077), .B(n3592), .C(n3628), .D(N8278), .Z(n2101) );
  CND3XL U12433 ( .A(n2102), .B(n2103), .C(n2104), .Z(N9324) );
  CANR2X1 U12434 ( .A(N2076), .B(n3592), .C(n3626), .D(N8279), .Z(n2104) );
  CND3XL U12435 ( .A(n3167), .B(n3168), .C(n3169), .Z(N10000) );
  CND3XL U12436 ( .A(n2132), .B(n2133), .C(n2134), .Z(N10345) );
  CANR2X1 U12437 ( .A(N3097), .B(n3594), .C(n3628), .D(N7258), .Z(n2134) );
  CND2X1 U12438 ( .A(N6179), .B(n3693), .Z(n2133) );
  CANR2X1 U12439 ( .A(mem_data1[1021]), .B(n3898), .C(N9301), .D(n3674), .Z(
        n2132) );
  CND3XL U12440 ( .A(n2135), .B(n2136), .C(n2137), .Z(N10344) );
  CANR2X1 U12441 ( .A(N3096), .B(n3594), .C(n3628), .D(N7259), .Z(n2137) );
  CND2X1 U12442 ( .A(N6178), .B(n3693), .Z(n2136) );
  CND3XL U12443 ( .A(n2138), .B(n2139), .C(n2140), .Z(N10343) );
  CANR2X1 U12444 ( .A(N3095), .B(n3594), .C(n3628), .D(N7260), .Z(n2140) );
  CND2X1 U12445 ( .A(N6177), .B(n3693), .Z(n2139) );
  CND3XL U12446 ( .A(n2141), .B(n2142), .C(n2143), .Z(N10342) );
  CANR2X1 U12447 ( .A(N3094), .B(n3594), .C(n3628), .D(N7261), .Z(n2143) );
  CND2X1 U12448 ( .A(N6176), .B(n3683), .Z(n2142) );
  CND3XL U12449 ( .A(n2144), .B(n2145), .C(n2146), .Z(N10341) );
  CANR2X1 U12450 ( .A(N3093), .B(n3594), .C(n3628), .D(N7262), .Z(n2146) );
  CND2X1 U12451 ( .A(N6175), .B(n3693), .Z(n2145) );
  CND3XL U12452 ( .A(n2147), .B(n2148), .C(n2149), .Z(N10340) );
  CANR2X1 U12453 ( .A(N3092), .B(n3594), .C(n3628), .D(N7263), .Z(n2149) );
  CND2X1 U12454 ( .A(N6174), .B(n3691), .Z(n2148) );
  CND3XL U12455 ( .A(n2150), .B(n2151), .C(n2152), .Z(N10339) );
  CANR2X1 U12456 ( .A(N3091), .B(n3594), .C(n3628), .D(N7264), .Z(n2152) );
  CND2X1 U12457 ( .A(N6173), .B(n3691), .Z(n2151) );
  CND3XL U12458 ( .A(n2153), .B(n2154), .C(n2155), .Z(N10338) );
  CANR2X1 U12459 ( .A(N3090), .B(n3594), .C(n3627), .D(N7265), .Z(n2155) );
  CND2X1 U12460 ( .A(N6172), .B(n3698), .Z(n2154) );
  CND3XL U12461 ( .A(n2156), .B(n2157), .C(n2158), .Z(N10337) );
  CANR2X1 U12462 ( .A(N3089), .B(n3594), .C(n3627), .D(N7266), .Z(n2158) );
  CND2X1 U12463 ( .A(N6171), .B(n3685), .Z(n2157) );
  CND3XL U12464 ( .A(n2159), .B(n2160), .C(n2161), .Z(N10336) );
  CANR2X1 U12465 ( .A(N3088), .B(n3593), .C(n3627), .D(N7267), .Z(n2161) );
  CND2X1 U12466 ( .A(N6170), .B(n3686), .Z(n2160) );
  CANR2X1 U12467 ( .A(mem_data1[1012]), .B(n3898), .C(N9292), .D(n3675), .Z(
        n2159) );
  CND3XL U12468 ( .A(n2162), .B(n2163), .C(n2164), .Z(N10335) );
  CANR2X1 U12469 ( .A(N3087), .B(n3593), .C(n3627), .D(N7268), .Z(n2164) );
  CND2X1 U12470 ( .A(N6169), .B(n3694), .Z(n2163) );
  CND3XL U12471 ( .A(n2165), .B(n2166), .C(n2167), .Z(N10334) );
  CANR2X1 U12472 ( .A(N3086), .B(n3593), .C(n3627), .D(N7269), .Z(n2167) );
  CND2X1 U12473 ( .A(N6168), .B(n3683), .Z(n2166) );
  CND3XL U12474 ( .A(n2168), .B(n2169), .C(n2170), .Z(N10333) );
  CANR2X1 U12475 ( .A(N3085), .B(n3593), .C(n3627), .D(N7270), .Z(n2170) );
  CND2X1 U12476 ( .A(N6167), .B(n3690), .Z(n2169) );
  CND3XL U12477 ( .A(n2171), .B(n2172), .C(n2173), .Z(N10332) );
  CANR2X1 U12478 ( .A(N3084), .B(n3593), .C(n3627), .D(N7271), .Z(n2173) );
  CND2X1 U12479 ( .A(N6166), .B(n3696), .Z(n2172) );
  CND3XL U12480 ( .A(n2174), .B(n2175), .C(n2176), .Z(N10331) );
  CND2X1 U12481 ( .A(N6165), .B(n3694), .Z(n2175) );
  CND3XL U12482 ( .A(n2177), .B(n2178), .C(n2179), .Z(N10330) );
  CND3XL U12483 ( .A(n2129), .B(n2130), .C(n2131), .Z(N10346) );
  CANR2X1 U12484 ( .A(N3098), .B(n3594), .C(n3628), .D(N7257), .Z(n2131) );
  CND2X1 U12485 ( .A(N6180), .B(n3693), .Z(n2130) );
  CND3XL U12486 ( .A(n2126), .B(n2127), .C(n2128), .Z(N10347) );
  CANR2X1 U12487 ( .A(N3099), .B(n3594), .C(n3628), .D(N7256), .Z(n2128) );
  CND2X1 U12488 ( .A(N6181), .B(n3693), .Z(n2127) );
  CAN2X1 U12489 ( .A(datain0[4]), .B(n4389), .Z(n5477) );
  CAN2X1 U12490 ( .A(datain0[3]), .B(n4389), .Z(n5473) );
  CAN2X1 U12491 ( .A(datain0[9]), .B(n4389), .Z(n5504) );
  CAN2X1 U12492 ( .A(datain0[7]), .B(n4389), .Z(n5492) );
  CAN2X1 U12493 ( .A(datain0[6]), .B(n4389), .Z(n5487) );
  CAN2X1 U12494 ( .A(datain0[11]), .B(n4388), .Z(n5516) );
  CAN2X1 U12495 ( .A(datain0[14]), .B(n4389), .Z(n5534) );
  CAN2X1 U12496 ( .A(datain0[13]), .B(n4389), .Z(n5528) );
  CAN2X1 U12497 ( .A(datain0[15]), .B(n4389), .Z(n5540) );
  CAN2X1 U12498 ( .A(datain0[18]), .B(n4389), .Z(n5560) );
  CAN2X1 U12499 ( .A(datain0[17]), .B(n4388), .Z(n5553) );
  CAN2X1 U12500 ( .A(datain0[16]), .B(n4389), .Z(n5546) );
  CAN2X1 U12501 ( .A(datain0[19]), .B(n4388), .Z(n5569) );
  CAN2X1 U12502 ( .A(datain0[26]), .B(n4388), .Z(n5618) );
  CAN2X1 U12503 ( .A(datain0[25]), .B(n4388), .Z(n5611) );
  CAN2X1 U12504 ( .A(datain0[5]), .B(n4389), .Z(n5482) );
  CAN2X1 U12505 ( .A(datain0[2]), .B(n4389), .Z(n5469) );
  CAN2X1 U12506 ( .A(datain0[0]), .B(n4389), .Z(n5464) );
  CAN2X1 U12507 ( .A(datain0[1]), .B(n4389), .Z(n5466) );
  CAN2X1 U12508 ( .A(datain0[8]), .B(n4389), .Z(n5497) );
  CAN2X1 U12509 ( .A(datain0[10]), .B(n4389), .Z(n5510) );
  CANR2X1 U12510 ( .A(N6222), .B(n3594), .C(N2066), .D(n3637), .Z(n2124) );
  CIVX2 U12511 ( .A(mem_data1[413]), .Z(n3743) );
  CNR2X1 U12512 ( .A(n4435), .B(pushin0), .Z(n73) );
  CNR2IX1 U12513 ( .B(mem_data1[1023]), .A(n3857), .Z(n6558) );
  CNR2X1 U12514 ( .A(lenout[0]), .B(lenout[1]), .Z(n15731) );
  CNR3XL U12515 ( .A(n52), .B(N10376), .C(n51), .Z(dataout[0]) );
  CNR2X1 U12516 ( .A(lenout[3]), .B(n15737), .Z(N10376) );
  CNR3XL U12517 ( .A(n52), .B(N10377), .C(n50), .Z(dataout[1]) );
  CNR2X1 U12518 ( .A(lenout[3]), .B(n15738), .Z(N10377) );
  CNR3XL U12519 ( .A(n52), .B(N10378), .C(n49), .Z(dataout[2]) );
  CNR2X1 U12520 ( .A(lenout[3]), .B(n15733), .Z(N10378) );
  CNR3XL U12521 ( .A(n52), .B(N10379), .C(n48), .Z(dataout[3]) );
  CNR2X1 U12522 ( .A(lenout[3]), .B(lenout[2]), .Z(N10379) );
  CNR3XL U12523 ( .A(n52), .B(N10380), .C(n47), .Z(dataout[4]) );
  CNR2X1 U12524 ( .A(n15734), .B(lenout[3]), .Z(N10380) );
  CNR3XL U12525 ( .A(n52), .B(N10381), .C(n46), .Z(dataout[5]) );
  CNR2X1 U12526 ( .A(n15735), .B(lenout[3]), .Z(N10381) );
  CNR3XL U12527 ( .A(n52), .B(N10382), .C(n45), .Z(dataout[6]) );
  CNR2X1 U12528 ( .A(n15736), .B(lenout[3]), .Z(N10382) );
  CNR3XL U12529 ( .A(n52), .B(n4438), .C(n44), .Z(dataout[7]) );
  CNR3XL U12530 ( .A(n52), .B(N10384), .C(n43), .Z(dataout[8]) );
  CND2X1 U12531 ( .A(n15737), .B(lenout[3]), .Z(N10384) );
  CNR3XL U12532 ( .A(n52), .B(N10385), .C(n42), .Z(dataout[9]) );
  CND2X1 U12533 ( .A(n15738), .B(lenout[3]), .Z(N10385) );
  CNR3XL U12534 ( .A(n52), .B(N10386), .C(n41), .Z(dataout[10]) );
  CND2X1 U12535 ( .A(n15733), .B(lenout[3]), .Z(N10386) );
  CNR3XL U12536 ( .A(n52), .B(N10387), .C(n40), .Z(dataout[11]) );
  CND2X1 U12537 ( .A(lenout[2]), .B(lenout[3]), .Z(N10387) );
  CNR3XL U12538 ( .A(n52), .B(N10388), .C(n39), .Z(dataout[12]) );
  CND2X1 U12539 ( .A(n15734), .B(lenout[3]), .Z(N10388) );
  CNR3XL U12540 ( .A(n52), .B(N10389), .C(n38), .Z(dataout[13]) );
  CND2X1 U12541 ( .A(n15735), .B(lenout[3]), .Z(N10389) );
  CNR3XL U12542 ( .A(n52), .B(N10390), .C(n37), .Z(dataout[14]) );
  CND2X1 U12543 ( .A(n15736), .B(lenout[3]), .Z(N10390) );
  CND2X1 U12544 ( .A(lenout[1]), .B(lenout[0]), .Z(n15732) );
  CIVX2 U12545 ( .A(rst), .Z(n4415) );
  CIVXL U12546 ( .A(n3534), .Z(n3270) );
  CIVXL U12547 ( .A(n3536), .Z(n3271) );
  CIVXL U12548 ( .A(n3538), .Z(n3272) );
  CIVXL U12549 ( .A(n3539), .Z(n3273) );
  CIVXL U12550 ( .A(n3540), .Z(n3274) );
  CIVXL U12551 ( .A(n3541), .Z(n3275) );
  CIVXL U12552 ( .A(n3542), .Z(n3276) );
  CIVXL U12553 ( .A(n3543), .Z(n3277) );
  CIVXL U12554 ( .A(n3543), .Z(n3278) );
  CIVXL U12555 ( .A(n3543), .Z(n3279) );
  CIVXL U12556 ( .A(n3543), .Z(n3280) );
  CIVXL U12557 ( .A(n3543), .Z(n3281) );
  CIVXL U12558 ( .A(n3543), .Z(n3282) );
  CIVXL U12559 ( .A(n3543), .Z(n3283) );
  CIVXL U12560 ( .A(n3543), .Z(n3284) );
  CIVXL U12561 ( .A(n3543), .Z(n3285) );
  CIVXL U12562 ( .A(n3544), .Z(n3286) );
  CIVXL U12563 ( .A(n3544), .Z(n3287) );
  CIVXL U12564 ( .A(n3544), .Z(n3288) );
  CIVXL U12565 ( .A(n3544), .Z(n3289) );
  CIVXL U12566 ( .A(n3544), .Z(n3290) );
  CIVXL U12567 ( .A(n3544), .Z(n3291) );
  CIVXL U12568 ( .A(n3544), .Z(n3292) );
  CIVXL U12569 ( .A(n3545), .Z(n3293) );
  CIVXL U12570 ( .A(n3545), .Z(n3294) );
  CIVXL U12571 ( .A(n3545), .Z(n3295) );
  CIVXL U12572 ( .A(n3545), .Z(n3296) );
  CIVXL U12573 ( .A(n3545), .Z(n3297) );
  CIVXL U12574 ( .A(n3545), .Z(n3298) );
  CIVXL U12575 ( .A(n3545), .Z(n3299) );
  CIVXL U12576 ( .A(n3545), .Z(n3300) );
  CIVXL U12577 ( .A(n3545), .Z(n3301) );
  CIVXL U12578 ( .A(n3546), .Z(n3302) );
  CIVXL U12579 ( .A(n3546), .Z(n3303) );
  CIVXL U12580 ( .A(n3546), .Z(n3304) );
  CIVXL U12581 ( .A(n3546), .Z(n3305) );
  CIVXL U12582 ( .A(n3546), .Z(n3306) );
  CIVXL U12583 ( .A(n3546), .Z(n3307) );
  CIVXL U12584 ( .A(n3546), .Z(n3308) );
  CIVXL U12585 ( .A(n3546), .Z(n3309) );
  CIVXL U12586 ( .A(n3546), .Z(n3310) );
  CIVXL U12587 ( .A(n3546), .Z(n3311) );
  CIVXL U12588 ( .A(n3547), .Z(n3312) );
  CIVXL U12589 ( .A(n3547), .Z(n3313) );
  CIVXL U12590 ( .A(n3547), .Z(n3314) );
  CIVXL U12591 ( .A(n3547), .Z(n3315) );
  CIVXL U12592 ( .A(n3547), .Z(n3316) );
  CIVXL U12593 ( .A(n3547), .Z(n3317) );
  CIVXL U12594 ( .A(n3547), .Z(n3318) );
  CIVXL U12595 ( .A(n3547), .Z(n3319) );
  CIVXL U12596 ( .A(n3547), .Z(n3320) );
  CIVXL U12597 ( .A(n3547), .Z(n3321) );
  CIVXL U12598 ( .A(n3548), .Z(n3322) );
  CIVXL U12599 ( .A(n3548), .Z(n3323) );
  CIVXL U12600 ( .A(n3548), .Z(n3324) );
  CIVXL U12601 ( .A(n3548), .Z(n3325) );
  CIVXL U12602 ( .A(n3548), .Z(n3326) );
  CIVXL U12603 ( .A(n3548), .Z(n3327) );
  CIVXL U12604 ( .A(n3548), .Z(n3328) );
  CIVXL U12605 ( .A(n3548), .Z(n3329) );
  CIVXL U12606 ( .A(n3548), .Z(n3330) );
  CIVXL U12607 ( .A(n3548), .Z(n3331) );
  CIVXL U12608 ( .A(n3549), .Z(n3332) );
  CIVXL U12609 ( .A(n3549), .Z(n3333) );
  CIVXL U12610 ( .A(n3549), .Z(n3334) );
  CIVXL U12611 ( .A(n3549), .Z(n3335) );
  CIVXL U12612 ( .A(n3549), .Z(n3336) );
  CIVXL U12613 ( .A(n3549), .Z(n3337) );
  CIVXL U12614 ( .A(n3549), .Z(n3338) );
  CIVXL U12615 ( .A(n3549), .Z(n3339) );
  CIVXL U12616 ( .A(n3549), .Z(n3340) );
  CIVXL U12617 ( .A(n3550), .Z(n3341) );
  CIVXL U12618 ( .A(n3550), .Z(n3342) );
  CIVXL U12619 ( .A(n3550), .Z(n3343) );
  CIVXL U12620 ( .A(n3550), .Z(n3344) );
  CIVXL U12621 ( .A(n3550), .Z(n3345) );
  CIVXL U12622 ( .A(n3550), .Z(n3346) );
  CIVXL U12623 ( .A(n3550), .Z(n3347) );
  CIVXL U12624 ( .A(n3550), .Z(n3348) );
  CIVXL U12625 ( .A(n3550), .Z(n3349) );
  CIVXL U12626 ( .A(n3550), .Z(n3350) );
  CIVXL U12627 ( .A(n3551), .Z(n3351) );
  CIVXL U12628 ( .A(n3551), .Z(n3352) );
  CIVXL U12629 ( .A(n3551), .Z(n3353) );
  CIVXL U12630 ( .A(n3551), .Z(n3354) );
  CIVXL U12631 ( .A(n3551), .Z(n3355) );
  CIVXL U12632 ( .A(n3551), .Z(n3356) );
  CIVXL U12633 ( .A(n3551), .Z(n3357) );
  CIVXL U12634 ( .A(n3551), .Z(n3358) );
  CIVXL U12635 ( .A(n3551), .Z(n3359) );
  CIVXL U12636 ( .A(n3551), .Z(n3360) );
  CIVXL U12637 ( .A(n3552), .Z(n3361) );
  CIVXL U12638 ( .A(n3552), .Z(n3362) );
  CIVXL U12639 ( .A(n3552), .Z(n3363) );
  CIVXL U12640 ( .A(n3552), .Z(n3364) );
  CIVXL U12641 ( .A(n3552), .Z(n3365) );
  CIVXL U12642 ( .A(n3552), .Z(n3366) );
  CIVXL U12643 ( .A(n3552), .Z(n3367) );
  CIVXL U12644 ( .A(n3552), .Z(n3368) );
  CIVXL U12645 ( .A(n3553), .Z(n3369) );
  CIVXL U12646 ( .A(n3553), .Z(n3370) );
  CIVXL U12647 ( .A(n3553), .Z(n3371) );
  CIVXL U12648 ( .A(n3553), .Z(n3372) );
  CIVXL U12649 ( .A(n3553), .Z(n3373) );
  CIVXL U12650 ( .A(n3553), .Z(n3374) );
  CIVXL U12651 ( .A(n3553), .Z(n3375) );
  CIVXL U12652 ( .A(n3553), .Z(n3376) );
  CIVXL U12653 ( .A(n3553), .Z(n3377) );
  CIVXL U12654 ( .A(n3553), .Z(n3378) );
  CIVXL U12655 ( .A(n3554), .Z(n3379) );
  CIVXL U12656 ( .A(n3554), .Z(n3380) );
  CIVXL U12657 ( .A(n3554), .Z(n3381) );
  CIVXL U12658 ( .A(n3554), .Z(n3382) );
  CIVXL U12659 ( .A(n3554), .Z(n3383) );
  CIVXL U12660 ( .A(n3554), .Z(n3384) );
  CIVXL U12661 ( .A(n3555), .Z(n3385) );
  CIVXL U12662 ( .A(n3555), .Z(n3386) );
  CIVXL U12663 ( .A(n3555), .Z(n3387) );
  CIVXL U12664 ( .A(n3555), .Z(n3388) );
  CIVXL U12665 ( .A(n3555), .Z(n3389) );
  CIVXL U12666 ( .A(n3555), .Z(n3390) );
  CIVXL U12667 ( .A(n3555), .Z(n3391) );
  CIVXL U12668 ( .A(n3555), .Z(n3392) );
  CIVXL U12669 ( .A(n3555), .Z(n3393) );
  CIVXL U12670 ( .A(n3555), .Z(n3394) );
  CIVXL U12671 ( .A(n3556), .Z(n3395) );
  CIVXL U12672 ( .A(n3556), .Z(n3396) );
  CIVXL U12673 ( .A(n3556), .Z(n3397) );
  CIVXL U12674 ( .A(n3556), .Z(n3398) );
  CIVXL U12675 ( .A(n3556), .Z(n3399) );
  CIVXL U12676 ( .A(n3556), .Z(n3400) );
  CIVXL U12677 ( .A(n3556), .Z(n3401) );
  CIVXL U12678 ( .A(n3556), .Z(n3402) );
  CIVXL U12679 ( .A(n3556), .Z(n3403) );
  CIVXL U12680 ( .A(n3556), .Z(n3404) );
  CIVXL U12681 ( .A(n3557), .Z(n3405) );
  CIVXL U12682 ( .A(n3557), .Z(n3406) );
  CIVXL U12683 ( .A(n3557), .Z(n3407) );
  CIVXL U12684 ( .A(n3557), .Z(n3408) );
  CIVXL U12685 ( .A(n3557), .Z(n3409) );
  CIVXL U12686 ( .A(n3557), .Z(n3410) );
  CIVXL U12687 ( .A(n3557), .Z(n3411) );
  CIVXL U12688 ( .A(n3557), .Z(n3412) );
  CIVXL U12689 ( .A(n3557), .Z(n3413) );
  CIVXL U12690 ( .A(n3557), .Z(n3414) );
  CIVXL U12691 ( .A(n3558), .Z(n3415) );
  CIVXL U12692 ( .A(n3558), .Z(n3416) );
  CIVXL U12693 ( .A(n3558), .Z(n3417) );
  CIVXL U12694 ( .A(n3558), .Z(n3418) );
  CIVXL U12695 ( .A(n3558), .Z(n3419) );
  CIVXL U12696 ( .A(n3558), .Z(n3420) );
  CIVXL U12697 ( .A(n3558), .Z(n3421) );
  CIVXL U12698 ( .A(n3558), .Z(n3422) );
  CIVXL U12699 ( .A(n3558), .Z(n3423) );
  CIVXL U12700 ( .A(n3558), .Z(n3424) );
  CIVXL U12701 ( .A(n3559), .Z(n3425) );
  CIVXL U12702 ( .A(n3559), .Z(n3426) );
  CIVXL U12703 ( .A(n3559), .Z(n3427) );
  CIVXL U12704 ( .A(n3559), .Z(n3428) );
  CIVXL U12705 ( .A(n3559), .Z(n3429) );
  CIVXL U12706 ( .A(n3559), .Z(n3430) );
  CIVXL U12707 ( .A(n3559), .Z(n3431) );
  CIVXL U12708 ( .A(n3559), .Z(n3432) );
  CIVXL U12709 ( .A(n3559), .Z(n3433) );
  CIVXL U12710 ( .A(n3559), .Z(n3434) );
  CIVXL U12711 ( .A(n3560), .Z(n3435) );
  CIVXL U12712 ( .A(n3560), .Z(n3436) );
  CIVXL U12713 ( .A(n3560), .Z(n3437) );
  CIVXL U12714 ( .A(n3560), .Z(n3438) );
  CIVXL U12715 ( .A(n3560), .Z(n3439) );
  CIVXL U12716 ( .A(n3560), .Z(n3440) );
  CIVXL U12717 ( .A(n3560), .Z(n3441) );
  CIVXL U12718 ( .A(n3560), .Z(n3442) );
  CIVXL U12719 ( .A(n3560), .Z(n3443) );
  CIVXL U12720 ( .A(n3560), .Z(n3444) );
  CIVXL U12721 ( .A(n3561), .Z(n3445) );
  CIVXL U12722 ( .A(n3561), .Z(n3446) );
  CIVXL U12723 ( .A(n3561), .Z(n3447) );
  CIVXL U12724 ( .A(n3561), .Z(n3448) );
  CIVXL U12725 ( .A(n3561), .Z(n3449) );
  CIVXL U12726 ( .A(n3561), .Z(n3450) );
  CIVXL U12727 ( .A(n3561), .Z(n3451) );
  CIVXL U12728 ( .A(n3561), .Z(n3452) );
  CIVXL U12729 ( .A(n3561), .Z(n3453) );
  CIVXL U12730 ( .A(n3561), .Z(n3454) );
  CIVXL U12731 ( .A(n3562), .Z(n3455) );
  CIVXL U12732 ( .A(n3562), .Z(n3456) );
  CIVXL U12733 ( .A(n3562), .Z(n3457) );
  CIVXL U12734 ( .A(n3562), .Z(n3458) );
  CIVXL U12735 ( .A(n3562), .Z(n3459) );
  CIVXL U12736 ( .A(n3562), .Z(n3460) );
  CIVXL U12737 ( .A(n3562), .Z(n3461) );
  CIVXL U12738 ( .A(n3562), .Z(n3462) );
  CIVXL U12739 ( .A(n3562), .Z(n3463) );
  CIVXL U12740 ( .A(n3562), .Z(n3464) );
  CIVXL U12741 ( .A(n3563), .Z(n3465) );
  CIVXL U12742 ( .A(n3563), .Z(n3466) );
  CIVXL U12743 ( .A(n3563), .Z(n3467) );
  CIVXL U12744 ( .A(n3563), .Z(n3468) );
  CIVXL U12745 ( .A(n3563), .Z(n3469) );
  CIVXL U12746 ( .A(n3563), .Z(n3470) );
  CIVXL U12747 ( .A(n3563), .Z(n3471) );
  CIVXL U12748 ( .A(n3563), .Z(n3472) );
  CIVXL U12749 ( .A(n3563), .Z(n3473) );
  CIVXL U12750 ( .A(n3563), .Z(n3474) );
  CIVXL U12751 ( .A(n3564), .Z(n3475) );
  CIVXL U12752 ( .A(n3564), .Z(n3476) );
  CIVXL U12753 ( .A(n3564), .Z(n3477) );
  CIVXL U12754 ( .A(n3564), .Z(n3478) );
  CIVXL U12755 ( .A(n3564), .Z(n3479) );
  CIVXL U12756 ( .A(n3564), .Z(n3480) );
  CIVXL U12757 ( .A(n3564), .Z(n3481) );
  CIVXL U12758 ( .A(n3564), .Z(n3482) );
  CIVXL U12759 ( .A(n3564), .Z(n3483) );
  CIVXL U12760 ( .A(n3564), .Z(n3484) );
  CIVXL U12761 ( .A(n3565), .Z(n3485) );
  CIVXL U12762 ( .A(n3565), .Z(n3486) );
  CIVXL U12763 ( .A(n3565), .Z(n3487) );
  CIVXL U12764 ( .A(n3565), .Z(n3488) );
  CIVXL U12765 ( .A(n3565), .Z(n3489) );
  CIVXL U12766 ( .A(n3565), .Z(n3490) );
  CIVXL U12767 ( .A(n3565), .Z(n3491) );
  CIVXL U12768 ( .A(n3565), .Z(n3492) );
  CIVXL U12769 ( .A(n3565), .Z(n3493) );
  CIVXL U12770 ( .A(n3565), .Z(n3494) );
  CIVXL U12771 ( .A(n3566), .Z(n3495) );
  CIVXL U12772 ( .A(n3566), .Z(n3496) );
  CIVXL U12773 ( .A(n3566), .Z(n3497) );
  CIVXL U12774 ( .A(n3566), .Z(n3498) );
  CIVXL U12775 ( .A(n3566), .Z(n3499) );
  CIVXL U12776 ( .A(n3566), .Z(n3500) );
  CIVXL U12777 ( .A(n3566), .Z(n3501) );
  CIVXL U12778 ( .A(n3566), .Z(n3502) );
  CIVXL U12779 ( .A(n3566), .Z(n3503) );
  CIVXL U12780 ( .A(n3566), .Z(n3504) );
  CIVXL U12781 ( .A(n3567), .Z(n3505) );
  CIVXL U12782 ( .A(n3567), .Z(n3506) );
  CIVXL U12783 ( .A(n3567), .Z(n3507) );
  CIVXL U12784 ( .A(n3567), .Z(n3508) );
  CIVXL U12785 ( .A(n3567), .Z(n3509) );
  CIVXL U12786 ( .A(n3567), .Z(n3510) );
  CIVXL U12787 ( .A(n3567), .Z(n3511) );
  CIVXL U12788 ( .A(n3567), .Z(n3512) );
  CIVXL U12789 ( .A(n3567), .Z(n3513) );
  CIVXL U12790 ( .A(n3567), .Z(n3514) );
  CIVXL U12791 ( .A(n3568), .Z(n3515) );
  CIVXL U12792 ( .A(n3568), .Z(n3516) );
  CIVXL U12793 ( .A(n3568), .Z(n3517) );
  CIVXL U12794 ( .A(n3568), .Z(n3518) );
  CIVXL U12795 ( .A(n3568), .Z(n3519) );
  CIVXL U12796 ( .A(n3568), .Z(n3520) );
  CIVXL U12797 ( .A(n3568), .Z(n3521) );
  CIVXL U12798 ( .A(n3568), .Z(n3522) );
  CIVXL U12799 ( .A(n3568), .Z(n3523) );
  CIVXL U12800 ( .A(n3568), .Z(n3524) );
  CIVXL U12801 ( .A(n3569), .Z(n3525) );
  CIVXL U12802 ( .A(n3569), .Z(n3526) );
  CIVXL U12803 ( .A(n3569), .Z(n3527) );
  CIVXL U12804 ( .A(n3569), .Z(n3528) );
  CIVXL U12805 ( .A(n3569), .Z(n3529) );
  CIVXL U12806 ( .A(n3569), .Z(n3530) );
  CIVXL U12807 ( .A(n3569), .Z(n3531) );
  CIVXL U12808 ( .A(n3569), .Z(n3532) );
  CIVX1 U12809 ( .A(n3897), .Z(n3534) );
  CIVX1 U12810 ( .A(n3897), .Z(n3535) );
  CIVX1 U12811 ( .A(n3897), .Z(n3536) );
  CIVX1 U12812 ( .A(n3897), .Z(n3537) );
  CIVX1 U12813 ( .A(n3897), .Z(n3538) );
  CIVX1 U12814 ( .A(n3897), .Z(n3539) );
  CIVX1 U12815 ( .A(n3897), .Z(n3540) );
  CIVX1 U12816 ( .A(n3897), .Z(n3541) );
  CIVX1 U12817 ( .A(n3897), .Z(n3542) );
  CIVX1 U12818 ( .A(n3897), .Z(n3543) );
  CIVX1 U12819 ( .A(n3897), .Z(n3544) );
  CIVX1 U12820 ( .A(n3897), .Z(n3545) );
  CIVX1 U12821 ( .A(n3897), .Z(n3546) );
  CIVX1 U12822 ( .A(n3897), .Z(n3547) );
  CIVX1 U12823 ( .A(n3897), .Z(n3548) );
  CIVX1 U12824 ( .A(n3897), .Z(n3549) );
  CIVX1 U12825 ( .A(n3897), .Z(n3550) );
  CIVX1 U12826 ( .A(n3897), .Z(n3551) );
  CIVX1 U12827 ( .A(n3897), .Z(n3552) );
  CIVX1 U12828 ( .A(n3897), .Z(n3553) );
  CIVX1 U12829 ( .A(n3897), .Z(n3554) );
  CIVX1 U12830 ( .A(n3897), .Z(n3555) );
  CIVX1 U12831 ( .A(n3897), .Z(n3556) );
  CIVX1 U12832 ( .A(n3897), .Z(n3557) );
  CIVX1 U12833 ( .A(n3897), .Z(n3558) );
  CIVX1 U12834 ( .A(n3897), .Z(n3559) );
  CIVX1 U12835 ( .A(n3897), .Z(n3560) );
  CIVX1 U12836 ( .A(n3897), .Z(n3561) );
  CIVX1 U12837 ( .A(n3897), .Z(n3562) );
  CIVX1 U12838 ( .A(n3897), .Z(n3563) );
  CIVX1 U12839 ( .A(n3897), .Z(n3564) );
  CIVX1 U12840 ( .A(n3897), .Z(n3565) );
  CIVX1 U12841 ( .A(n3897), .Z(n3566) );
  CIVX1 U12842 ( .A(n3897), .Z(n3567) );
  CIVX1 U12843 ( .A(n3897), .Z(n3568) );
  CIVX1 U12844 ( .A(n3897), .Z(n3569) );
  CMXI2X1 U12845 ( .A0(n13316), .A1(n13322), .S(n3750), .Z(n13329) );
  CND3XL U12846 ( .A(n1226), .B(n1227), .C(n1228), .Z(N9616) );
  CND3XL U12847 ( .A(n1220), .B(n1221), .C(n1222), .Z(N9618) );
  CND3XL U12848 ( .A(n896), .B(n897), .C(n898), .Z(N9726) );
  CANR2X1 U12849 ( .A(mem_data1[402]), .B(n3898), .C(N8682), .D(n3681), .Z(
        n896) );
  CMXI2X1 U12850 ( .A0(n13328), .A1(n13337), .S(n3750), .Z(n13344) );
  CND3XL U12851 ( .A(n1223), .B(n1224), .C(n1225), .Z(N9617) );
  CND3XL U12852 ( .A(n1193), .B(n1194), .C(n1195), .Z(N9627) );
  CND3XL U12853 ( .A(n1187), .B(n1188), .C(n1189), .Z(N9629) );
  CND3XL U12854 ( .A(n1160), .B(n1161), .C(n1162), .Z(N9638) );
  CND3XL U12855 ( .A(n1154), .B(n1155), .C(n1156), .Z(N9640) );
  CND3XL U12856 ( .A(n854), .B(n855), .C(n856), .Z(N9740) );
  CANR2X1 U12857 ( .A(mem_data1[408]), .B(n3898), .C(n3678), .D(N8688), .Z(
        n878) );
  CANR2X1 U12858 ( .A(mem_data1[404]), .B(n3898), .C(n3678), .D(N8684), .Z(
        n890) );
  CMX2XL U12859 ( .A0(n4757), .A1(n4756), .S(n3203), .Z(n4879) );
  CND2X1 U12860 ( .A(n4819), .B(n3740), .Z(n4930) );
  CND3XL U12861 ( .A(n1232), .B(n1233), .C(n1234), .Z(N9614) );
  CEOX1 U12862 ( .A(N135), .B(mem_data1[117]), .Z(N8162) );
  CND2X1 U12863 ( .A(n3728), .B(n4879), .Z(n6225) );
  CND2X1 U12864 ( .A(n4879), .B(n3739), .Z(n6008) );
  CANR2X1 U12865 ( .A(mem_data1[440]), .B(n3898), .C(n3678), .D(N8720), .Z(
        n782) );
  CEOX1 U12866 ( .A(N377), .B(mem_data1[359]), .Z(N7920) );
  CMXI2X1 U12867 ( .A0(n13750), .A1(n13756), .S(n3750), .Z(n13763) );
  CMXI2X1 U12868 ( .A0(n13413), .A1(n13419), .S(n3750), .Z(n13426) );
  CMXI2X1 U12869 ( .A0(n13756), .A1(n13762), .S(n3750), .Z(n13769) );
  CND3XL U12870 ( .A(n1004), .B(n1005), .C(n1006), .Z(N9690) );
  CANR2X1 U12871 ( .A(mem_data1[374]), .B(n3898), .C(n3678), .D(N8654), .Z(
        n980) );
  CND2X1 U12872 ( .A(n3764), .B(n4227), .Z(n3747) );
  CANR2X1 U12873 ( .A(N2427), .B(n3604), .C(n3637), .D(N7928), .Z(n1051) );
  CND2X1 U12874 ( .A(n3728), .B(n4900), .Z(n5112) );
  CND2X1 U12875 ( .A(n4900), .B(n3731), .Z(n6397) );
  CND3XL U12876 ( .A(n1364), .B(n1365), .C(n1366), .Z(N9570) );
  CND3XL U12877 ( .A(n767), .B(n768), .C(n769), .Z(N9769) );
  CANR2X1 U12878 ( .A(mem_data1[245]), .B(n3898), .C(N8525), .D(n3682), .Z(
        n1367) );
  CANR2X1 U12879 ( .A(N2432), .B(n3604), .C(n3637), .D(N7923), .Z(n1036) );
  CEOX1 U12880 ( .A(N374), .B(mem_data1[356]), .Z(N7923) );
  CND3XL U12881 ( .A(n629), .B(n630), .C(n631), .Z(N9815) );
  CND3XL U12882 ( .A(n623), .B(n624), .C(n625), .Z(N9817) );
  CEOX1 U12883 ( .A(N511), .B(mem_data1[493]), .Z(N7786) );
  CANR2X1 U12884 ( .A(N2363), .B(n3604), .C(n3637), .D(N7992), .Z(n1243) );
  CANR2XL U12885 ( .A(N2390), .B(n3604), .C(n3638), .D(N7965), .Z(n1162) );
  CMXI2XL U12886 ( .A0(n4663), .A1(n4666), .S(n4223), .Z(n3699) );
  CMXI2XL U12887 ( .A0(n4663), .A1(n4666), .S(n4221), .Z(n4702) );
  CANR2XL U12888 ( .A(N2392), .B(n3604), .C(n3638), .D(N7963), .Z(n1156) );
  CEOX1 U12889 ( .A(N120), .B(mem_data1[102]), .Z(N8177) );
  CANR2X1 U12890 ( .A(mem_data1[98]), .B(n3898), .C(N8378), .D(n3679), .Z(
        n1808) );
  CANR2X1 U12891 ( .A(mem_data1[90]), .B(n3898), .C(N8370), .D(n3679), .Z(
        n1832) );
  CND3XL U12892 ( .A(n887), .B(n888), .C(n889), .Z(N9729) );
  CND3XL U12893 ( .A(n626), .B(n627), .C(n628), .Z(N9816) );
  CEOX1 U12894 ( .A(N510), .B(mem_data1[492]), .Z(N7787) );
  CND2X1 U12895 ( .A(N5509), .B(n3695), .Z(n1050) );
  CMXI2X1 U12896 ( .A0(n13407), .A1(n13413), .S(n3750), .Z(n13420) );
  CANR2X1 U12897 ( .A(mem_data1[415]), .B(n3898), .C(n3678), .D(N8695), .Z(
        n857) );
  CANR2X1 U12898 ( .A(mem_data1[407]), .B(n3898), .C(n3678), .D(N8687), .Z(
        n881) );
  CND2X1 U12899 ( .A(N5514), .B(n3698), .Z(n1035) );
  CANR2X1 U12900 ( .A(N2122), .B(n3604), .C(n3637), .D(N8233), .Z(n1966) );
  CANR2X1 U12901 ( .A(mem_data1[439]), .B(n3898), .C(n3678), .D(N8719), .Z(
        n785) );
  CANR2X1 U12902 ( .A(mem_data1[435]), .B(n3898), .C(n3678), .D(N8715), .Z(
        n797) );
  CND2X1 U12903 ( .A(N5513), .B(n3698), .Z(n1038) );
  CMXI2XL U12904 ( .A0(n4675), .A1(n4673), .S(n3892), .Z(n3700) );
  CMXI2XL U12905 ( .A0(n4675), .A1(n4673), .S(n3892), .Z(n4711) );
  CANR2X1 U12906 ( .A(N2386), .B(n3604), .C(n3638), .D(N7969), .Z(n1174) );
  CMXI2X1 U12907 ( .A0(n13765), .A1(n13771), .S(n3750), .Z(n13781) );
  CANR2X1 U12908 ( .A(mem_data1[434]), .B(n3898), .C(n3678), .D(N8714), .Z(
        n800) );
  CANR2X1 U12909 ( .A(mem_data1[436]), .B(n3898), .C(n3678), .D(N8716), .Z(
        n794) );
  CANR2X1 U12910 ( .A(mem_data1[442]), .B(n3898), .C(n3679), .D(N8722), .Z(
        n776) );
  CANR2X1 U12911 ( .A(mem_data1[444]), .B(n3898), .C(n3679), .D(N8724), .Z(
        n770) );
  CANR2X1 U12912 ( .A(N2238), .B(n3604), .C(n3637), .D(N8117), .Z(n1618) );
  CND2X1 U12913 ( .A(n4810), .B(n3200), .Z(n4911) );
  CMXI2X1 U12914 ( .A0(n14175), .A1(n13907), .S(n3534), .Z(N8324) );
  CANR2X1 U12915 ( .A(N2250), .B(n3604), .C(n3637), .D(N8105), .Z(n1582) );
  CIVX2 U12916 ( .A(n4295), .Z(n4238) );
  CIVX2 U12917 ( .A(n4295), .Z(n4237) );
  CANR2X1 U12918 ( .A(N2572), .B(n3604), .C(n3637), .D(N7783), .Z(n616) );
  CMX2XL U12919 ( .A0(N7783), .A1(N7782), .S(n4252), .Z(n10948) );
  CEOX1 U12920 ( .A(N514), .B(mem_data1[496]), .Z(N7783) );
  CANR2X1 U12921 ( .A(N2314), .B(n3604), .C(n3638), .D(N8041), .Z(n1390) );
  CMX2XL U12922 ( .A0(N8042), .A1(N8041), .S(n4244), .Z(n10079) );
  CEOX1 U12923 ( .A(N256), .B(mem_data1[238]), .Z(N8041) );
  CANR2X1 U12924 ( .A(mem_data1[370]), .B(n3898), .C(n3678), .D(N8650), .Z(
        n992) );
  CANR2X1 U12925 ( .A(mem_data1[378]), .B(n3898), .C(n3678), .D(N8658), .Z(
        n968) );
  CANR2X1 U12926 ( .A(N2575), .B(n3604), .C(n3637), .D(N7780), .Z(n607) );
  CMX2XL U12927 ( .A0(N7780), .A1(N7779), .S(n4252), .Z(n10957) );
  CMX2XL U12928 ( .A0(N7781), .A1(N7780), .S(n4252), .Z(n10954) );
  CEOX1 U12929 ( .A(N517), .B(mem_data1[499]), .Z(N7780) );
  CND3XL U12930 ( .A(n764), .B(n765), .C(n766), .Z(N9770) );
  CANR2X1 U12931 ( .A(mem_data1[438]), .B(n3898), .C(n3678), .D(N8718), .Z(
        n788) );
  CMXI2X1 U12932 ( .A0(n13901), .A1(n13877), .S(n3534), .Z(N8720) );
  CANR2X1 U12933 ( .A(N2185), .B(n3604), .C(n3637), .D(N8170), .Z(n1777) );
  CMX2XL U12934 ( .A0(N8171), .A1(N8170), .S(n4287), .Z(n9652) );
  CEOX1 U12935 ( .A(N127), .B(mem_data1[109]), .Z(N8170) );
  CND3XL U12936 ( .A(n851), .B(n852), .C(n853), .Z(N9741) );
  CND3XL U12937 ( .A(n2090), .B(n2091), .C(n2092), .Z(N9328) );
  CIVXL U12938 ( .A(n4685), .Z(n3702) );
  CND2X1 U12939 ( .A(n3765), .B(n3891), .Z(n3703) );
  CMXI2X1 U12940 ( .A0(n13679), .A1(n13652), .S(n3535), .Z(N8654) );
  CANR2XL U12941 ( .A(N2389), .B(n3604), .C(n3638), .D(N7966), .Z(n1165) );
  CND2X1 U12942 ( .A(n5219), .B(n3204), .Z(n5320) );
  CMXI2X1 U12943 ( .A0(n13846), .A1(n13852), .S(n3750), .Z(n3704) );
  CMXI2X1 U12944 ( .A0(n13854), .A1(n13880), .S(n3343), .Z(N8713) );
  CEOX1 U12945 ( .A(N372), .B(mem_data1[354]), .Z(N7925) );
  CEOX1 U12946 ( .A(N392), .B(mem_data1[374]), .Z(N7905) );
  CEOX1 U12947 ( .A(N264), .B(mem_data1[246]), .Z(N8033) );
  CMXI2X1 U12948 ( .A0(n13394), .A1(n13410), .S(n3750), .Z(n13417) );
  CANR2X1 U12949 ( .A(N2266), .B(n3604), .C(n3637), .D(N8089), .Z(n1534) );
  CEOX1 U12950 ( .A(N380), .B(mem_data1[362]), .Z(N7917) );
  CMX2X1 U12951 ( .A0(n5206), .A1(n5308), .S(n3729), .Z(n3705) );
  CND3XL U12952 ( .A(n1157), .B(n1158), .C(n1159), .Z(N9639) );
  CND3XL U12953 ( .A(n1151), .B(n1152), .C(n1153), .Z(N9641) );
  CND3XL U12954 ( .A(n806), .B(n807), .C(n808), .Z(N9756) );
  CMXI2X1 U12955 ( .A0(n13845), .A1(n13868), .S(n3343), .Z(N8710) );
  CMXI2XL U12956 ( .A0(n4687), .A1(n4685), .S(n3891), .Z(n3706) );
  CMXI2XL U12957 ( .A0(n3701), .A1(n4687), .S(n3765), .Z(n4719) );
  CMXI2X1 U12958 ( .A0(n5024), .A1(n5123), .S(n3761), .Z(n3712) );
  CANR2XL U12959 ( .A(N2391), .B(n3604), .C(n3638), .D(N7964), .Z(n1159) );
  CANR2X1 U12960 ( .A(N2372), .B(n3604), .C(n3637), .D(N7983), .Z(n1216) );
  CANR2X1 U12961 ( .A(N2515), .B(n3604), .C(n3637), .D(N7840), .Z(n787) );
  CANR2X1 U12962 ( .A(N2111), .B(n3604), .C(n3637), .D(N8244), .Z(n1999) );
  CANR2X1 U12963 ( .A(mem_data1[33]), .B(n3898), .C(N8313), .D(n3679), .Z(
        n2003) );
  CMX2XL U12964 ( .A0(N8245), .A1(N8244), .S(n4246), .Z(n10094) );
  CMX2XL U12965 ( .A0(N8244), .A1(N8243), .S(n4245), .Z(n10127) );
  CMXI2X1 U12966 ( .A0(n13910), .A1(n13883), .S(n3535), .Z(N8722) );
  CMXI2X1 U12967 ( .A0(n13916), .A1(n13889), .S(n3535), .Z(N8724) );
  CANR2X1 U12968 ( .A(N2555), .B(n3604), .C(n3638), .D(N7800), .Z(n667) );
  CANR2X1 U12969 ( .A(mem_data1[363]), .B(n3898), .C(N8643), .D(n3680), .Z(
        n1013) );
  CANR2X1 U12970 ( .A(mem_data1[365]), .B(n3898), .C(N8645), .D(n3680), .Z(
        n1007) );
  CMXI2X1 U12971 ( .A0(n13691), .A1(n13664), .S(n3535), .Z(N8658) );
  CMX2X1 U12972 ( .A0(N7832), .A1(N7831), .S(n3862), .Z(n3707) );
  CANR2X1 U12973 ( .A(N2177), .B(n3604), .C(n3637), .D(N8178), .Z(n1801) );
  CMX2XL U12974 ( .A0(N8179), .A1(N8178), .S(n4286), .Z(n12237) );
  CEOX1 U12975 ( .A(N119), .B(mem_data1[101]), .Z(N8178) );
  CANR2X1 U12976 ( .A(mem_data1[339]), .B(n3898), .C(n3679), .D(N8619), .Z(
        n1085) );
  CANR2X1 U12977 ( .A(mem_data1[341]), .B(n3898), .C(n3678), .D(N8621), .Z(
        n1079) );
  CMXI2X1 U12978 ( .A0(n13614), .A1(n13620), .S(n3750), .Z(n13627) );
  CMX2X1 U12979 ( .A0(n5354), .A1(n5253), .S(n3735), .Z(n5426) );
  CANR2X1 U12980 ( .A(N2239), .B(n3604), .C(n3637), .D(N8116), .Z(n1615) );
  CMX2XL U12981 ( .A0(N8117), .A1(N8116), .S(n4280), .Z(n9825) );
  CMX2XL U12982 ( .A0(N8116), .A1(N8115), .S(n4280), .Z(n9828) );
  CANR2X1 U12983 ( .A(mem_data1[340]), .B(n3898), .C(n3678), .D(N8620), .Z(
        n1082) );
  CANR2X1 U12984 ( .A(mem_data1[342]), .B(n3898), .C(n3678), .D(N8622), .Z(
        n1076) );
  CMXI2X1 U12985 ( .A0(n13623), .A1(n13617), .S(n4180), .Z(n3708) );
  CND2X1 U12986 ( .A(n5209), .B(n3214), .Z(n5312) );
  CND3XL U12987 ( .A(n863), .B(n864), .C(n865), .Z(N9737) );
  CANR2X1 U12988 ( .A(N2303), .B(n3604), .C(n3638), .D(N8052), .Z(n1423) );
  CMX2XL U12989 ( .A0(N8052), .A1(N8051), .S(n4245), .Z(n10046) );
  CMX2XL U12990 ( .A0(N8053), .A1(N8052), .S(n4245), .Z(n10043) );
  CEOX1 U12991 ( .A(N245), .B(mem_data1[227]), .Z(N8052) );
  CANR2XL U12992 ( .A(N2234), .B(n3605), .C(n3638), .D(N8121), .Z(n1630) );
  CANR2X1 U12993 ( .A(mem_data1[156]), .B(n3898), .C(N8436), .D(n3681), .Z(
        n1634) );
  CANR2XL U12994 ( .A(N2507), .B(n3605), .C(n3638), .D(N7848), .Z(n811) );
  CND2X1 U12995 ( .A(n5223), .B(n3204), .Z(n5324) );
  CND2X1 U12996 ( .A(n5157), .B(n3207), .Z(n5224) );
  CMXI2X1 U12997 ( .A0(n13843), .A1(n13849), .S(n3750), .Z(n13856) );
  CANR2X1 U12998 ( .A(N2451), .B(n3604), .C(n3637), .D(N7904), .Z(n979) );
  CEOX1 U12999 ( .A(N393), .B(mem_data1[375]), .Z(N7904) );
  CANR2X1 U13000 ( .A(N2175), .B(n3604), .C(n3637), .D(N8180), .Z(n1807) );
  CMX2XL U13001 ( .A0(N8180), .A1(N8179), .S(n3878), .Z(n12270) );
  CMX2XL U13002 ( .A0(N8181), .A1(N8180), .S(n3879), .Z(n12236) );
  CEOX1 U13003 ( .A(N117), .B(mem_data1[99]), .Z(N8180) );
  CANR2X1 U13004 ( .A(mem_data1[345]), .B(n3898), .C(n3678), .D(N8625), .Z(
        n1067) );
  CANR2X1 U13005 ( .A(mem_data1[353]), .B(n3898), .C(n3678), .D(N8633), .Z(
        n1043) );
  CANR2X1 U13006 ( .A(mem_data1[343]), .B(n3898), .C(n3678), .D(N8623), .Z(
        n1073) );
  CMX2X1 U13007 ( .A0(n5350), .A1(n5249), .S(n3735), .Z(n5424) );
  CANR2X1 U13008 ( .A(n3898), .B(mem_data1[4]), .C(N8284), .D(n3680), .Z(n2090) );
  CIVXL U13009 ( .A(n14073), .Z(n4424) );
  CND2X1 U13010 ( .A(n5161), .B(n3203), .Z(n5228) );
  CANR2X1 U13011 ( .A(mem_data1[346]), .B(n3898), .C(n3678), .D(N8626), .Z(
        n1064) );
  CANR2X1 U13012 ( .A(mem_data1[354]), .B(n3898), .C(n3678), .D(N8634), .Z(
        n1040) );
  CMXI2X1 U13013 ( .A0(n13770), .A1(n13746), .S(n3536), .Z(N8680) );
  CANR2X1 U13014 ( .A(N2192), .B(n3604), .C(n3638), .D(N8163), .Z(n1756) );
  CMX2XL U13015 ( .A0(N8163), .A1(N8162), .S(n4286), .Z(n9665) );
  CEOX1 U13016 ( .A(N134), .B(mem_data1[116]), .Z(N8163) );
  CANR2X1 U13017 ( .A(mem_data1[344]), .B(n3898), .C(n3678), .D(N8624), .Z(
        n1070) );
  CMXI2X1 U13018 ( .A0(n13533), .A1(n13542), .S(n3750), .Z(n13549) );
  CANR2XL U13019 ( .A(N2190), .B(n3605), .C(n3639), .D(N8165), .Z(n1762) );
  CEOX1 U13020 ( .A(N132), .B(mem_data1[114]), .Z(N8165) );
  CEOX1 U13021 ( .A(N144), .B(mem_data1[126]), .Z(N8153) );
  CMX2XL U13022 ( .A0(N7976), .A1(N7975), .S(n4240), .Z(n10298) );
  CANR2X1 U13023 ( .A(N2379), .B(n3604), .C(n3637), .D(N7976), .Z(n1195) );
  CMXI2X1 U13024 ( .A0(n13539), .A1(n13545), .S(n3750), .Z(n13552) );
  CANR2XL U13025 ( .A(N2501), .B(n3604), .C(n3638), .D(N7854), .Z(n829) );
  CANR2XL U13026 ( .A(N2388), .B(n3604), .C(n3638), .D(N7967), .Z(n1168) );
  CMX2XL U13027 ( .A0(N7968), .A1(N7967), .S(n4239), .Z(n10322) );
  CANR2XL U13028 ( .A(N2520), .B(n3605), .C(n3638), .D(N7835), .Z(n772) );
  CANR2X1 U13029 ( .A(mem_data1[58]), .B(n3898), .C(N8338), .D(n3679), .Z(
        n1928) );
  CANR2X1 U13030 ( .A(mem_data1[489]), .B(n3898), .C(N8769), .D(n3680), .Z(
        n635) );
  CANR2X1 U13031 ( .A(N2500), .B(n3604), .C(n3637), .D(N7855), .Z(n832) );
  CND2X1 U13032 ( .A(n3727), .B(n5263), .Z(n5365) );
  CANR2X1 U13033 ( .A(N2431), .B(n3604), .C(n3637), .D(N7924), .Z(n1039) );
  CMX2XL U13034 ( .A0(N7924), .A1(N7923), .S(n4261), .Z(n10476) );
  CEOX1 U13035 ( .A(N373), .B(mem_data1[355]), .Z(N7924) );
  CMXI2X1 U13036 ( .A0(n13971), .A1(n14037), .S(n3750), .Z(n14108) );
  CANR2X1 U13037 ( .A(mem_data1[488]), .B(n3898), .C(N8768), .D(n3681), .Z(
        n638) );
  CANR2XL U13038 ( .A(N2560), .B(n3605), .C(n3639), .D(N7795), .Z(n652) );
  CEOX1 U13039 ( .A(mem_data1[484]), .B(N502), .Z(N7795) );
  CANR2XL U13040 ( .A(N2496), .B(n3604), .C(n3638), .D(N7859), .Z(n844) );
  CANR2X1 U13041 ( .A(mem_data1[490]), .B(n3898), .C(N8770), .D(n3681), .Z(
        n632) );
  CANR2X1 U13042 ( .A(N2198), .B(n3604), .C(n3637), .D(N8157), .Z(n1738) );
  CMXI2X1 U13043 ( .A0(n13995), .A1(n14001), .S(n3750), .Z(n14011) );
  CANR2XL U13044 ( .A(N2195), .B(n3605), .C(n3639), .D(N8160), .Z(n1747) );
  CANR2X1 U13045 ( .A(mem_data1[361]), .B(n3898), .C(N8641), .D(n3680), .Z(
        n1019) );
  CANR2XL U13046 ( .A(N2367), .B(n3605), .C(n3638), .D(N7988), .Z(n1231) );
  CAN2X1 U13047 ( .A(n4790), .B(n3203), .Z(n4856) );
  CANR2X1 U13048 ( .A(mem_data1[116]), .B(n3898), .C(N8396), .D(n3680), .Z(
        n1754) );
  CMXI2XL U13049 ( .A0(n13563), .A1(n13572), .S(n3750), .Z(n3709) );
  CANR2X1 U13050 ( .A(mem_data1[362]), .B(n3898), .C(N8642), .D(n3680), .Z(
        n1016) );
  CANR2XL U13051 ( .A(N2495), .B(n3605), .C(n3638), .D(N7860), .Z(n847) );
  CMXI2X1 U13052 ( .A0(n13998), .A1(n14007), .S(n3750), .Z(n14014) );
  CMXI2XL U13053 ( .A0(n4583), .A1(n4586), .S(n3194), .Z(n3710) );
  CMXI2XL U13054 ( .A0(n4583), .A1(n4586), .S(n3188), .Z(n4515) );
  CANR2X1 U13055 ( .A(mem_data1[119]), .B(n3898), .C(N8399), .D(n3680), .Z(
        n1745) );
  CANR2XL U13056 ( .A(N2407), .B(n3604), .C(n3638), .D(N7948), .Z(n1111) );
  CMX2XL U13057 ( .A0(N7948), .A1(N7947), .S(n4229), .Z(n10395) );
  CMX2XL U13058 ( .A0(N7949), .A1(N7948), .S(n4280), .Z(n10392) );
  CMXI2X1 U13059 ( .A0(n13563), .A1(n13572), .S(n3750), .Z(n13579) );
  CMXI2X1 U13060 ( .A0(n12763), .A1(n12769), .S(lenin0[1]), .Z(n12776) );
  CANR2X1 U13061 ( .A(N2323), .B(n3604), .C(n3638), .D(N8032), .Z(n1363) );
  CANR2XL U13062 ( .A(N2384), .B(n3605), .C(n3638), .D(N7971), .Z(n1180) );
  CANR2X1 U13063 ( .A(mem_data1[493]), .B(n3898), .C(N8773), .D(n3681), .Z(
        n623) );
  CMXI2XL U13064 ( .A0(n12760), .A1(n12751), .S(n4199), .Z(n3711) );
  CMXI2XL U13065 ( .A0(n12760), .A1(n12751), .S(n4199), .Z(n12767) );
  CANR2XL U13066 ( .A(N2513), .B(n3605), .C(n3638), .D(N7842), .Z(n793) );
  CMX2XL U13067 ( .A0(N7975), .A1(N7974), .S(n4239), .Z(n10301) );
  CANR2X1 U13068 ( .A(N2381), .B(n3604), .C(n3637), .D(N7974), .Z(n1189) );
  CANR2XL U13069 ( .A(n3691), .B(N8265), .C(mem_data1[14]), .D(n3250), .Z(n56)
         );
  CANR2X1 U13070 ( .A(N2090), .B(n3604), .C(n3637), .D(N8265), .Z(n2062) );
  CND2X1 U13071 ( .A(n4888), .B(n3735), .Z(n6203) );
  CND2X1 U13072 ( .A(n3723), .B(n4888), .Z(n4784) );
  CANR2XL U13073 ( .A(N2517), .B(n3605), .C(n3638), .D(N7838), .Z(n781) );
  CANR2X1 U13074 ( .A(mem_data1[441]), .B(n3898), .C(n3679), .D(N8721), .Z(
        n779) );
  CANR2X1 U13075 ( .A(mem_data1[437]), .B(n3898), .C(n3678), .D(N8717), .Z(
        n791) );
  CANR2XL U13076 ( .A(N2476), .B(n3605), .C(n3638), .D(N7879), .Z(n904) );
  CANR2X1 U13077 ( .A(mem_data1[398]), .B(n3898), .C(N8678), .D(n3681), .Z(
        n908) );
  CANR2X1 U13078 ( .A(N6230), .B(n2105), .C(n3898), .D(n4386), .Z(n2109) );
  CNR2X1 U13079 ( .A(n5113), .B(n3896), .Z(n5141) );
  CNR2IX1 U13080 ( .B(datain0[31]), .A(n4386), .Z(n5090) );
  CNR2IX1 U13081 ( .B(datain0[29]), .A(n4386), .Z(n5076) );
  CNR2IX1 U13082 ( .B(datain0[30]), .A(n4386), .Z(n5083) );
  CNR2IX1 U13083 ( .B(datain0[27]), .A(n4386), .Z(n5062) );
  CNR2IX1 U13084 ( .B(datain0[25]), .A(n4386), .Z(n5048) );
  CNR2IX1 U13085 ( .B(datain0[28]), .A(n4386), .Z(n5069) );
  CNR2IX1 U13086 ( .B(datain0[26]), .A(n4386), .Z(n5055) );
  CANR2XL U13087 ( .A(N2374), .B(n3605), .C(n3638), .D(N7981), .Z(n1210) );
  CMXI2X1 U13088 ( .A0(n14001), .A1(n14010), .S(n3750), .Z(n14017) );
  CANR2XL U13089 ( .A(N2429), .B(n3604), .C(n3638), .D(N7926), .Z(n1045) );
  CMX2XL U13090 ( .A0(N7927), .A1(N7926), .S(n4237), .Z(n10467) );
  CEOX1 U13091 ( .A(N371), .B(mem_data1[353]), .Z(N7926) );
  CMXI2X1 U13092 ( .A0(n13334), .A1(n13340), .S(n3750), .Z(n13347) );
  CMXI2X1 U13093 ( .A0(n12798), .A1(n12774), .S(n3536), .Z(N8394) );
  CMXI2X1 U13094 ( .A0(n12804), .A1(n12780), .S(n3537), .Z(N8396) );
  CEOX1 U13095 ( .A(N263), .B(mem_data1[245]), .Z(N8034) );
  CANR2X1 U13096 ( .A(mem_data1[230]), .B(n3898), .C(N8510), .D(n3680), .Z(
        n1412) );
  CMXI2X1 U13097 ( .A0(n13819), .A1(n13825), .S(n3750), .Z(n13832) );
  CANR2X1 U13098 ( .A(mem_data1[243]), .B(n3898), .C(N8523), .D(n3680), .Z(
        n1373) );
  CMXI2X1 U13099 ( .A0(n13246), .A1(n13219), .S(n3537), .Z(N8525) );
  CMXI2X1 U13100 ( .A0(n13831), .A1(n13837), .S(n3750), .Z(n13847) );
  CEOX1 U13101 ( .A(N270), .B(mem_data1[252]), .Z(N8027) );
  CMXI2X1 U13102 ( .A0(n14007), .A1(n14013), .S(n3750), .Z(n14020) );
  CMXI2X1 U13103 ( .A0(n13169), .A1(n13175), .S(n3750), .Z(n13182) );
  CANR2X1 U13104 ( .A(N2347), .B(n3604), .C(n3638), .D(N8008), .Z(n1291) );
  CMX2XL U13105 ( .A0(N8008), .A1(N8007), .S(n4228), .Z(n10190) );
  CANR2XL U13106 ( .A(N2394), .B(n3604), .C(n3638), .D(N7961), .Z(n1150) );
  CMXI2X1 U13107 ( .A0(n13172), .A1(n13178), .S(n3750), .Z(n13185) );
  CANR2XL U13108 ( .A(N2170), .B(n3605), .C(n3639), .D(N8185), .Z(n1822) );
  CMX2XL U13109 ( .A0(N8185), .A1(N8184), .S(n3868), .Z(n12104) );
  CMX2XL U13110 ( .A0(N8186), .A1(N8185), .S(n3881), .Z(n12071) );
  CEOX1 U13111 ( .A(N112), .B(mem_data1[94]), .Z(N8185) );
  CANR2XL U13112 ( .A(N2491), .B(n3605), .C(n3638), .D(N7864), .Z(n859) );
  CMX2XL U13113 ( .A0(N7864), .A1(N7863), .S(n4256), .Z(n10681) );
  CMX2XL U13114 ( .A0(N7865), .A1(N7864), .S(n4256), .Z(n10678) );
  CEOX1 U13115 ( .A(N265), .B(mem_data1[247]), .Z(N8032) );
  CEOX1 U13116 ( .A(N272), .B(mem_data1[254]), .Z(N8025) );
  CANR2XL U13117 ( .A(N2458), .B(n3605), .C(n3638), .D(N7897), .Z(n958) );
  CANR2XL U13118 ( .A(N2298), .B(n3605), .C(n3638), .D(N8057), .Z(n1438) );
  CMX2XL U13119 ( .A0(N8058), .A1(N8057), .S(n4246), .Z(n10025) );
  CANR2XL U13120 ( .A(N2365), .B(n3605), .C(n3638), .D(N7990), .Z(n1237) );
  CMX2XL U13121 ( .A0(N7991), .A1(N7990), .S(n4240), .Z(n10247) );
  CANR2XL U13122 ( .A(N2376), .B(n3605), .C(n3638), .D(N7979), .Z(n1204) );
  CMX2XL U13123 ( .A0(N7979), .A1(N7978), .S(n4240), .Z(n10286) );
  CND2X1 U13124 ( .A(N5444), .B(n3696), .Z(n1245) );
  CND2X1 U13125 ( .A(n5201), .B(n3208), .Z(n5303) );
  CANR2X1 U13126 ( .A(mem_data1[250]), .B(n3898), .C(N8530), .D(n3682), .Z(
        n1352) );
  CANR2XL U13127 ( .A(N2411), .B(n3604), .C(n3638), .D(N7944), .Z(n1099) );
  CMX2XL U13128 ( .A0(N7944), .A1(N7943), .S(n4238), .Z(n10410) );
  CMX2XL U13129 ( .A0(N7945), .A1(N7944), .S(n4238), .Z(n10407) );
  CANR2XL U13130 ( .A(N2378), .B(n3605), .C(n3638), .D(N7977), .Z(n1198) );
  CMX2XL U13131 ( .A0(N7978), .A1(N7977), .S(n4240), .Z(n10289) );
  CMX2XL U13132 ( .A0(N7977), .A1(N7976), .S(n4240), .Z(n10295) );
  CMX2XL U13133 ( .A0(N7849), .A1(N7848), .S(n4231), .Z(n10729) );
  CMX2XL U13134 ( .A0(N7850), .A1(N7849), .S(n4235), .Z(n10726) );
  CANR2X1 U13135 ( .A(N2506), .B(n3604), .C(n3637), .D(N7849), .Z(n814) );
  CANR2XL U13136 ( .A(N2373), .B(n3605), .C(n3638), .D(N7982), .Z(n1213) );
  CANR2X1 U13137 ( .A(mem_data1[251]), .B(n3898), .C(N8531), .D(n3682), .Z(
        n1349) );
  CND3XL U13138 ( .A(n959), .B(n960), .C(n961), .Z(N9705) );
  CANR2XL U13139 ( .A(N2351), .B(n3605), .C(n3638), .D(N8004), .Z(n1279) );
  CMX2XL U13140 ( .A0(N8004), .A1(N8003), .S(n4241), .Z(n10205) );
  CMX2XL U13141 ( .A0(N8005), .A1(N8004), .S(n4241), .Z(n10202) );
  CANR2XL U13142 ( .A(N2557), .B(n3605), .C(n3639), .D(N7798), .Z(n661) );
  CMX2XL U13143 ( .A0(N7799), .A1(N7798), .S(n4280), .Z(n10894) );
  CEOX1 U13144 ( .A(mem_data1[481]), .B(N499), .Z(N7798) );
  CANR2X1 U13145 ( .A(mem_data1[350]), .B(n3898), .C(n3678), .D(N8630), .Z(
        n1052) );
  CANR2XL U13146 ( .A(N2504), .B(n3604), .C(n3638), .D(N7851), .Z(n820) );
  CMX2XL U13147 ( .A0(N7851), .A1(N7850), .S(n4253), .Z(n10723) );
  CANR2X1 U13148 ( .A(mem_data1[359]), .B(n3898), .C(n3678), .D(N8639), .Z(
        n1025) );
  CANR2X1 U13149 ( .A(mem_data1[348]), .B(n3898), .C(n3678), .D(N8628), .Z(
        n1058) );
  CMX2X1 U13150 ( .A0(n5198), .A1(n5299), .S(n3729), .Z(n3713) );
  CND2X1 U13151 ( .A(n5197), .B(n3214), .Z(n5299) );
  CANR2XL U13152 ( .A(N2522), .B(n3605), .C(n3638), .D(N7833), .Z(n766) );
  CMXI2X1 U13153 ( .A0(n13613), .A1(n13586), .S(n3538), .Z(N8634) );
  CANR2XL U13154 ( .A(N2502), .B(n3604), .C(n3638), .D(N7853), .Z(n826) );
  CMX2XL U13155 ( .A0(N7853), .A1(N7852), .S(n4253), .Z(n10717) );
  CND3XL U13156 ( .A(n962), .B(n963), .C(n964), .Z(N9704) );
  CANR2X1 U13157 ( .A(mem_data1[349]), .B(n3898), .C(n3678), .D(N8629), .Z(
        n1055) );
  CEOX1 U13158 ( .A(N267), .B(mem_data1[249]), .Z(N8030) );
  CANR2X1 U13159 ( .A(mem_data1[242]), .B(n3898), .C(N8522), .D(n3679), .Z(
        n1376) );
  CANR2X1 U13160 ( .A(mem_data1[234]), .B(n3898), .C(N8514), .D(n3680), .Z(
        n1400) );
  CANR2X1 U13161 ( .A(mem_data1[252]), .B(n3898), .C(N8532), .D(n3682), .Z(
        n1346) );
  CANR2XL U13162 ( .A(N2559), .B(n3605), .C(n3639), .D(N7796), .Z(n655) );
  CMX2XL U13163 ( .A0(N7796), .A1(N7795), .S(n4235), .Z(n10906) );
  CEOX1 U13164 ( .A(N501), .B(mem_data1[483]), .Z(N7796) );
  CANR2XL U13165 ( .A(N2385), .B(n3605), .C(n3638), .D(N7970), .Z(n1177) );
  CMX2XL U13166 ( .A0(N7971), .A1(N7970), .S(n4239), .Z(n10313) );
  CMX2XL U13167 ( .A0(N7970), .A1(N7969), .S(n4239), .Z(n10316) );
  CANR2XL U13168 ( .A(N2518), .B(n3605), .C(n3638), .D(N7837), .Z(n778) );
  CMXI2X1 U13169 ( .A0(n13181), .A1(n13187), .S(n3750), .Z(n13194) );
  CANR2XL U13170 ( .A(N2415), .B(n3604), .C(n3638), .D(N7940), .Z(n1087) );
  CMX2XL U13171 ( .A0(N7940), .A1(N7939), .S(n4238), .Z(n10422) );
  CMX2XL U13172 ( .A0(N7941), .A1(N7940), .S(n4238), .Z(n10419) );
  CMXI2X1 U13173 ( .A0(n13917), .A1(n13923), .S(n3750), .Z(n13930) );
  CMXI2X1 U13174 ( .A0(n13226), .A1(n13235), .S(n3750), .Z(n13242) );
  CMXI2X1 U13175 ( .A0(n13610), .A1(n13583), .S(n3538), .Z(N8633) );
  CMXI2X1 U13176 ( .A0(n13262), .A1(n13271), .S(n3750), .Z(n13278) );
  CMX2XL U13177 ( .A0(N7966), .A1(N7965), .S(n4239), .Z(n10338) );
  CMX2XL U13178 ( .A0(N7967), .A1(N7966), .S(n4239), .Z(n10335) );
  CANR2X1 U13179 ( .A(mem_data1[253]), .B(n3898), .C(N8533), .D(n3681), .Z(
        n1343) );
  CANR2XL U13180 ( .A(N2305), .B(n3605), .C(n3638), .D(N8050), .Z(n1417) );
  CMX2XL U13181 ( .A0(N8051), .A1(N8050), .S(n4245), .Z(n10049) );
  CMXI2XL U13182 ( .A0(n4603), .A1(n4602), .S(n3194), .Z(n4638) );
  CMX2XL U13183 ( .A0(N7964), .A1(N7963), .S(n4254), .Z(n10344) );
  CMX2XL U13184 ( .A0(N7965), .A1(N7964), .S(n4234), .Z(n10341) );
  CANR2X1 U13185 ( .A(N2194), .B(n3604), .C(n3638), .D(N8161), .Z(n1750) );
  CMX2XL U13186 ( .A0(N8161), .A1(N8160), .S(n4286), .Z(n9673) );
  CMX2XL U13187 ( .A0(N8162), .A1(N8161), .S(n4286), .Z(n9669) );
  CEOX1 U13188 ( .A(N136), .B(mem_data1[118]), .Z(N8161) );
  CND2X1 U13189 ( .A(n5182), .B(n3207), .Z(n5249) );
  CANR2XL U13190 ( .A(N2516), .B(n3605), .C(n3638), .D(N7839), .Z(n784) );
  CMX2XL U13191 ( .A0(N7840), .A1(N7839), .S(n4231), .Z(n10759) );
  CMXI2X1 U13192 ( .A0(n3716), .A1(n5073), .S(n3765), .Z(n5145) );
  CMXI2X1 U13193 ( .A0(n13628), .A1(n13601), .S(n3539), .Z(N8639) );
  CANR2XL U13194 ( .A(N2343), .B(n3605), .C(n3638), .D(N8012), .Z(n1303) );
  CMX2XL U13195 ( .A0(N8012), .A1(N8011), .S(n4229), .Z(n10178) );
  CMX2XL U13196 ( .A0(N8013), .A1(N8012), .S(n4242), .Z(n10175) );
  CMXI2X1 U13197 ( .A0(n13482), .A1(n13488), .S(n3750), .Z(n13495) );
  CANR2X1 U13198 ( .A(mem_data1[469]), .B(n3898), .C(n3677), .D(N8749), .Z(
        n695) );
  CANR2X1 U13199 ( .A(mem_data1[473]), .B(n3898), .C(n3678), .D(N8753), .Z(
        n683) );
  CMX2XL U13200 ( .A0(N7852), .A1(N7851), .S(n4254), .Z(n10720) );
  CANR2X1 U13201 ( .A(N2503), .B(n3604), .C(n3637), .D(N7852), .Z(n823) );
  CND2X1 U13202 ( .A(n5203), .B(n3208), .Z(n5306) );
  CND2X1 U13203 ( .A(n5263), .B(n3735), .Z(n5436) );
  CMXI2X1 U13204 ( .A0(n13521), .A1(n13527), .S(n3750), .Z(n13534) );
  CMXI2X1 U13205 ( .A0(n13950), .A1(n13956), .S(n3750), .Z(n13963) );
  CANR2X1 U13206 ( .A(mem_data1[256]), .B(n3898), .C(N8536), .D(n3681), .Z(
        n1334) );
  CND3XL U13207 ( .A(n1049), .B(n1050), .C(n1051), .Z(N9675) );
  CMX2XL U13208 ( .A0(N7848), .A1(N7847), .S(n4232), .Z(n10732) );
  CANR2XL U13209 ( .A(N2173), .B(n3605), .C(n3639), .D(N8182), .Z(n1813) );
  CMX2XL U13210 ( .A0(N8183), .A1(N8182), .S(n3869), .Z(n12170) );
  CMX2XL U13211 ( .A0(N8182), .A1(N8181), .S(n3866), .Z(n12203) );
  CND2X1 U13212 ( .A(n4808), .B(n3202), .Z(n4909) );
  CANR2XL U13213 ( .A(N2514), .B(n3605), .C(n3639), .D(N7841), .Z(n790) );
  CMX2XL U13214 ( .A0(N7841), .A1(N7840), .S(n4232), .Z(n10756) );
  CANR2XL U13215 ( .A(N2519), .B(n3605), .C(n3639), .D(N7836), .Z(n775) );
  CMX2XL U13216 ( .A0(N7837), .A1(N7836), .S(n4232), .Z(n10771) );
  CND3XL U13217 ( .A(n1046), .B(n1047), .C(n1048), .Z(N9676) );
  CANR2XL U13218 ( .A(N2512), .B(n3605), .C(n3639), .D(N7843), .Z(n796) );
  CANR2X1 U13219 ( .A(mem_data1[257]), .B(n3898), .C(N8537), .D(n3681), .Z(
        n1331) );
  CMXI2XL U13220 ( .A0(n5094), .A1(n5037), .S(n4221), .Z(n3715) );
  CMXI2XL U13221 ( .A0(n5094), .A1(n5037), .S(n4226), .Z(n5130) );
  CMX2XL U13222 ( .A0(N7860), .A1(N7859), .S(n4252), .Z(n10693) );
  CANR2XL U13223 ( .A(N2186), .B(n3605), .C(n3639), .D(N8169), .Z(n1774) );
  CMX2XL U13224 ( .A0(N8170), .A1(N8169), .S(n4286), .Z(n9659) );
  CMX2XL U13225 ( .A0(N8169), .A1(N8168), .S(n4287), .Z(n9653) );
  CEOX1 U13226 ( .A(N128), .B(mem_data1[110]), .Z(N8169) );
  CANR2X1 U13227 ( .A(mem_data1[957]), .B(n3898), .C(N9237), .D(n3682), .Z(
        n2324) );
  CNR2X1 U13228 ( .A(n3840), .B(n6463), .Z(N849) );
  CNR2X1 U13229 ( .A(n3833), .B(n6463), .Z(N977) );
  CNR2X1 U13230 ( .A(n3763), .B(n6147), .Z(n6190) );
  CNR2IX1 U13231 ( .B(datain0[8]), .A(n4388), .Z(n4935) );
  CNR2IX1 U13232 ( .B(datain0[3]), .A(n4388), .Z(n6037) );
  CNR2IX1 U13233 ( .B(datain0[4]), .A(n4389), .Z(n6041) );
  CNR2IX1 U13234 ( .B(datain0[5]), .A(n4386), .Z(n6046) );
  CNR2IX1 U13235 ( .B(datain0[6]), .A(n4387), .Z(n6051) );
  CNR2IX1 U13236 ( .B(datain0[2]), .A(n4388), .Z(n6032) );
  CNR2IX1 U13237 ( .B(datain0[1]), .A(n4387), .Z(n6029) );
  CNR2IX1 U13238 ( .B(datain0[0]), .A(n4386), .Z(n6027) );
  CANR2X1 U13239 ( .A(mem_data1[320]), .B(n3898), .C(N8600), .D(n3679), .Z(
        n1142) );
  CANR2XL U13240 ( .A(N2371), .B(n3605), .C(n3638), .D(N7984), .Z(n1219) );
  CMX2XL U13241 ( .A0(N7984), .A1(N7983), .S(n4240), .Z(n10271) );
  CANR2XL U13242 ( .A(N2306), .B(n3605), .C(n3638), .D(N8049), .Z(n1414) );
  CANR2X1 U13243 ( .A(mem_data1[220]), .B(n3898), .C(N8500), .D(n3682), .Z(
        n1442) );
  CMX2XL U13244 ( .A0(N8050), .A1(N8049), .S(n4245), .Z(n10052) );
  CANR2XL U13245 ( .A(N2452), .B(n3605), .C(n3638), .D(N7903), .Z(n976) );
  CMX2XL U13246 ( .A0(N7904), .A1(N7903), .S(n4260), .Z(n10542) );
  CEOX1 U13247 ( .A(N394), .B(mem_data1[376]), .Z(N7903) );
  CIVX2 U13248 ( .A(n5181), .Z(n3716) );
  CIVXL U13249 ( .A(n5118), .Z(n3717) );
  CND2X1 U13250 ( .A(n3765), .B(n3891), .Z(n3718) );
  CND3XL U13251 ( .A(n1028), .B(n1029), .C(n1030), .Z(N9682) );
  CND2X1 U13252 ( .A(n6246), .B(n3735), .Z(n6348) );
  CNR2IX1 U13253 ( .B(n6178), .A(n3211), .Z(n6246) );
  CMXI2XL U13254 ( .A0(n4533), .A1(n6133), .S(n3764), .Z(n6178) );
  CANR2XL U13255 ( .A(N2475), .B(n3605), .C(n3638), .D(N7880), .Z(n907) );
  CANR2X1 U13256 ( .A(mem_data1[396]), .B(n3898), .C(N8676), .D(n3681), .Z(
        n914) );
  CMX2XL U13257 ( .A0(N7881), .A1(N7880), .S(n4258), .Z(n10617) );
  CMX2XL U13258 ( .A0(N7880), .A1(N7879), .S(n4257), .Z(n10620) );
  CANR2XL U13259 ( .A(N2449), .B(n3605), .C(n3638), .D(N7906), .Z(n985) );
  CEOX1 U13260 ( .A(N391), .B(mem_data1[373]), .Z(N7906) );
  CANR2XL U13261 ( .A(N2493), .B(n3605), .C(n3639), .D(N7862), .Z(n853) );
  CMX2XL U13262 ( .A0(N7863), .A1(N7862), .S(n4256), .Z(n10684) );
  CND3XL U13263 ( .A(n1034), .B(n1035), .C(n1036), .Z(N9680) );
  CANR2X1 U13264 ( .A(mem_data1[397]), .B(n3898), .C(N8677), .D(n3681), .Z(
        n911) );
  CANR2XL U13265 ( .A(N2471), .B(n3605), .C(n3638), .D(N7884), .Z(n919) );
  CANR2X1 U13266 ( .A(mem_data1[395]), .B(n3898), .C(N8675), .D(n3681), .Z(
        n917) );
  CMX2XL U13267 ( .A0(N7885), .A1(N7884), .S(n4258), .Z(n10605) );
  CMX2XL U13268 ( .A0(N7884), .A1(N7883), .S(n4258), .Z(n10608) );
  CND3XL U13269 ( .A(n1031), .B(n1032), .C(n1033), .Z(N9681) );
  CMXI2XL U13270 ( .A0(n5073), .A1(n5118), .S(n3891), .Z(n3719) );
  CANR2X1 U13271 ( .A(mem_data1[393]), .B(n3898), .C(N8673), .D(n3681), .Z(
        n923) );
  CANR2XL U13272 ( .A(N2567), .B(n3605), .C(n3638), .D(N7788), .Z(n631) );
  CMX2X1 U13273 ( .A0(N7789), .A1(N7788), .S(n3869), .Z(n13998) );
  CNIVX1 U13274 ( .A(n3721), .Z(n3722) );
  CNIVX1 U13275 ( .A(n3721), .Z(n3723) );
  CNIVX1 U13276 ( .A(n3721), .Z(n3724) );
  CNIVX1 U13277 ( .A(n3721), .Z(n3725) );
  CNIVX1 U13278 ( .A(wr_ptr[6]), .Z(n3726) );
  CNIVX1 U13279 ( .A(wr_ptr[6]), .Z(n3727) );
  CNIVX1 U13280 ( .A(wr_ptr[6]), .Z(n3728) );
  CNIVX1 U13281 ( .A(wr_ptr[6]), .Z(n3729) );
  CNIVX1 U13282 ( .A(wr_ptr[6]), .Z(n3730) );
  CNIVX1 U13283 ( .A(n3720), .Z(n3731) );
  CNIVX1 U13284 ( .A(n3720), .Z(n3732) );
  CNIVX1 U13285 ( .A(n3720), .Z(n3733) );
  CNIVX1 U13286 ( .A(n3720), .Z(n3734) );
  CNIVX1 U13287 ( .A(n3720), .Z(n3735) );
  CNIVX1 U13288 ( .A(n3720), .Z(n3736) );
  CNIVX1 U13289 ( .A(n3720), .Z(n3737) );
  CNIVX1 U13290 ( .A(n3720), .Z(n3738) );
  CNIVX1 U13291 ( .A(n3720), .Z(n3739) );
  CNIVX1 U13292 ( .A(n3720), .Z(n3740) );
  CANR2XL U13293 ( .A(N2319), .B(n3605), .C(n3638), .D(N8036), .Z(n1375) );
  CMX2X1 U13294 ( .A0(N8036), .A1(N8035), .S(n3875), .Z(n13172) );
  CNR2X1 U13295 ( .A(n3763), .B(n4227), .Z(n3741) );
  CIVX2 U13296 ( .A(n3754), .Z(n4227) );
  CANR2X1 U13297 ( .A(mem_data1[460]), .B(n3898), .C(N8740), .D(n3681), .Z(
        n722) );
  CANR2XL U13298 ( .A(N2440), .B(n3605), .C(n3638), .D(N7915), .Z(n1012) );
  CEOX1 U13299 ( .A(N382), .B(mem_data1[364]), .Z(N7915) );
  CND2X1 U13300 ( .A(n3722), .B(n5285), .Z(n5388) );
  CND2X1 U13301 ( .A(n5180), .B(n3201), .Z(n5247) );
  CND2X1 U13302 ( .A(n5285), .B(n3738), .Z(n5458) );
  CANR2XL U13303 ( .A(N2539), .B(n3605), .C(n3639), .D(N7816), .Z(n715) );
  CMX2XL U13304 ( .A0(N7816), .A1(N7815), .S(n4254), .Z(n10840) );
  CMX2XL U13305 ( .A0(N7817), .A1(N7816), .S(n4254), .Z(n10837) );
  CMXI2X1 U13306 ( .A0(n5066), .A1(n5114), .S(n3891), .Z(n5142) );
  CMXI2X1 U13307 ( .A0(n13914), .A1(n13920), .S(n3750), .Z(n13927) );
  CMXI2XL U13308 ( .A0(n4995), .A1(n5052), .S(n3891), .Z(n3742) );
  CMXI2XL U13309 ( .A0(n4995), .A1(n5052), .S(n3741), .Z(n5105) );
  CANR2XL U13310 ( .A(N2383), .B(n3605), .C(n3638), .D(N7972), .Z(n1183) );
  CMX2XL U13311 ( .A0(N7972), .A1(N7971), .S(n4239), .Z(n10310) );
  CANR2X1 U13312 ( .A(mem_data1[457]), .B(n3898), .C(N8737), .D(n3680), .Z(
        n731) );
  CMX2XL U13313 ( .A0(N7854), .A1(N7853), .S(n4255), .Z(n10714) );
  CMX2XL U13314 ( .A0(N7855), .A1(N7854), .S(n4254), .Z(n10711) );
  CND3XL U13315 ( .A(n1037), .B(n1038), .C(n1039), .Z(N9679) );
  CANR2XL U13316 ( .A(N2320), .B(n3605), .C(n3638), .D(N8035), .Z(n1372) );
  CEOX1 U13317 ( .A(N262), .B(mem_data1[244]), .Z(N8035) );
  CMXI2X1 U13318 ( .A0(n13324), .A1(n13297), .S(n3539), .Z(N8549) );
  CANR2X1 U13319 ( .A(mem_data1[461]), .B(n3898), .C(N8741), .D(n3680), .Z(
        n719) );
  CANR2XL U13320 ( .A(N2566), .B(n3605), .C(n3638), .D(N7789), .Z(n634) );
  CEOX1 U13321 ( .A(N508), .B(mem_data1[490]), .Z(N7789) );
  CMXI2X1 U13322 ( .A0(n13890), .A1(n13896), .S(n3750), .Z(n13903) );
  CANR2XL U13323 ( .A(N2453), .B(n3605), .C(n3638), .D(N7902), .Z(n973) );
  CMX2XL U13324 ( .A0(N7903), .A1(N7902), .S(n4260), .Z(n10545) );
  CEOX1 U13325 ( .A(N395), .B(mem_data1[377]), .Z(N7902) );
  CANR2X1 U13326 ( .A(mem_data1[277]), .B(n3898), .C(N8557), .D(n3679), .Z(
        n1271) );
  CANR2XL U13327 ( .A(N2479), .B(n3605), .C(n3638), .D(N7876), .Z(n895) );
  CANR2X1 U13328 ( .A(mem_data1[401]), .B(n3898), .C(N8681), .D(n3681), .Z(
        n899) );
  CMX2XL U13329 ( .A0(N7877), .A1(N7876), .S(n4257), .Z(n10632) );
  CMX2XL U13330 ( .A0(N7876), .A1(N7875), .S(n4257), .Z(n10635) );
  CANR2XL U13331 ( .A(N2442), .B(n3605), .C(n3638), .D(N7913), .Z(n1006) );
  CEOX1 U13332 ( .A(N384), .B(mem_data1[366]), .Z(N7913) );
  CMXI2X1 U13333 ( .A0(n5052), .A1(n5104), .S(n3891), .Z(n5136) );
  CANR2XL U13334 ( .A(N2455), .B(n3605), .C(n3638), .D(N7900), .Z(n967) );
  CANR2X1 U13335 ( .A(mem_data1[373]), .B(n3898), .C(n3678), .D(N8653), .Z(
        n983) );
  CANR2X1 U13336 ( .A(mem_data1[295]), .B(n3898), .C(n3678), .D(N8575), .Z(
        n1217) );
  CANR2X1 U13337 ( .A(mem_data1[299]), .B(n3898), .C(n3678), .D(N8579), .Z(
        n1205) );
  CANR2XL U13338 ( .A(N2437), .B(n3605), .C(n3638), .D(N7918), .Z(n1021) );
  CEOX1 U13339 ( .A(N379), .B(mem_data1[361]), .Z(N7918) );
  CMX2XL U13340 ( .A0(N7838), .A1(N7837), .S(n4233), .Z(n10765) );
  CMX2XL U13341 ( .A0(N7839), .A1(N7838), .S(n4229), .Z(n10762) );
  CANR2X1 U13342 ( .A(mem_data1[464]), .B(n3898), .C(N8744), .D(n3679), .Z(
        n710) );
  CMX2XL U13343 ( .A0(N7842), .A1(N7841), .S(n4234), .Z(n10753) );
  CMX2XL U13344 ( .A0(N7843), .A1(N7842), .S(n4233), .Z(n10750) );
  CMXI2X1 U13345 ( .A0(n13370), .A1(n13376), .S(n3750), .Z(n13383) );
  CENX1 U13346 ( .A(N431), .B(n3743), .Z(N7866) );
  CANR2X1 U13347 ( .A(mem_data1[309]), .B(n3898), .C(n3678), .D(N8589), .Z(
        n1175) );
  CANR2X1 U13348 ( .A(mem_data1[313]), .B(n3898), .C(n3678), .D(N8593), .Z(
        n1163) );
  CANR2X1 U13349 ( .A(mem_data1[273]), .B(n3898), .C(N8553), .D(n3679), .Z(
        n1283) );
  CANR2X1 U13350 ( .A(mem_data1[465]), .B(n3898), .C(N8745), .D(n3680), .Z(
        n707) );
  CANR2XL U13351 ( .A(N2450), .B(n3605), .C(n3638), .D(N7905), .Z(n982) );
  CMX2XL U13352 ( .A0(N7906), .A1(N7905), .S(n4260), .Z(n10536) );
  CMX2XL U13353 ( .A0(N7905), .A1(N7904), .S(n4260), .Z(n10539) );
  CMX2XL U13354 ( .A0(N7982), .A1(N7981), .S(n4240), .Z(n10277) );
  CMX2XL U13355 ( .A0(N7983), .A1(N7982), .S(n4240), .Z(n10274) );
  CANR2X1 U13356 ( .A(mem_data1[271]), .B(n3898), .C(N8551), .D(n3679), .Z(
        n1289) );
  CANR2XL U13357 ( .A(N2477), .B(n3605), .C(n3638), .D(N7878), .Z(n901) );
  CANR2X1 U13358 ( .A(mem_data1[399]), .B(n3898), .C(N8679), .D(n3681), .Z(
        n905) );
  CMX2XL U13359 ( .A0(N7879), .A1(N7878), .S(n4257), .Z(n10623) );
  CMX2XL U13360 ( .A0(N7878), .A1(N7877), .S(n4257), .Z(n10626) );
  CMXI2X1 U13361 ( .A0(n13416), .A1(n13422), .S(n3750), .Z(n13429) );
  CANR2X1 U13362 ( .A(mem_data1[385]), .B(n3898), .C(n3678), .D(N8665), .Z(
        n947) );
  CANR2X1 U13363 ( .A(mem_data1[377]), .B(n3898), .C(n3678), .D(N8657), .Z(
        n971) );
  CMXI2X1 U13364 ( .A0(n13653), .A1(n13659), .S(n3750), .Z(n13666) );
  CANR2XL U13365 ( .A(N2326), .B(n3605), .C(n3638), .D(N8029), .Z(n1354) );
  CANR2X1 U13366 ( .A(mem_data1[248]), .B(n3898), .C(N8528), .D(n3681), .Z(
        n1358) );
  CEOX1 U13367 ( .A(N268), .B(mem_data1[250]), .Z(N8029) );
  CANR2X1 U13368 ( .A(mem_data1[337]), .B(n3898), .C(N8617), .D(n3680), .Z(
        n1091) );
  CANR2XL U13369 ( .A(N2565), .B(n3605), .C(n3638), .D(N7790), .Z(n637) );
  CMX2XL U13370 ( .A0(N7790), .A1(N7789), .S(n4234), .Z(n10924) );
  CEOX1 U13371 ( .A(N507), .B(mem_data1[489]), .Z(N7790) );
  CANR2XL U13372 ( .A(N2315), .B(n3605), .C(n3638), .D(N8040), .Z(n1387) );
  CMX2XL U13373 ( .A0(N8040), .A1(N8039), .S(n4244), .Z(n10085) );
  CMX2XL U13374 ( .A0(N8041), .A1(N8040), .S(n4244), .Z(n10082) );
  CEOX1 U13375 ( .A(N257), .B(mem_data1[239]), .Z(N8040) );
  CANR2X1 U13376 ( .A(mem_data1[335]), .B(n3898), .C(N8615), .D(n3680), .Z(
        n1097) );
  CANR2XL U13377 ( .A(N2541), .B(n3605), .C(n3639), .D(N7814), .Z(n709) );
  CANR2X1 U13378 ( .A(mem_data1[463]), .B(n3898), .C(N8743), .D(n3680), .Z(
        n713) );
  CMX2XL U13379 ( .A0(N7815), .A1(N7814), .S(n4254), .Z(n10843) );
  CMX2XL U13380 ( .A0(N7814), .A1(N7813), .S(n4254), .Z(n10846) );
  CMX2XL U13381 ( .A0(N7836), .A1(N7835), .S(n4234), .Z(n10774) );
  CND3XL U13382 ( .A(n965), .B(n966), .C(n967), .Z(N9703) );
  CEOX1 U13383 ( .A(N397), .B(mem_data1[379]), .Z(N7900) );
  CANR2XL U13384 ( .A(N2322), .B(n3605), .C(n3638), .D(N8033), .Z(n1366) );
  CMX2XL U13385 ( .A0(N8033), .A1(N8032), .S(n4243), .Z(n10109) );
  CANR2X1 U13386 ( .A(mem_data1[409]), .B(n3898), .C(n3678), .D(N8689), .Z(
        n875) );
  CANR2X1 U13387 ( .A(mem_data1[278]), .B(n3898), .C(N8558), .D(n3679), .Z(
        n1268) );
  CANR2XL U13388 ( .A(N2456), .B(n3605), .C(n3638), .D(N7899), .Z(n964) );
  CMX2XL U13389 ( .A0(N7900), .A1(N7899), .S(n4259), .Z(n10554) );
  CEOX1 U13390 ( .A(N398), .B(mem_data1[380]), .Z(N7899) );
  CAN2XL U13391 ( .A(\r347/carry [4]), .B(n3757), .Z(\r347/carry [5]) );
  CNR2XL U13392 ( .A(n5747), .B(n3757), .Z(n5813) );
  CNR2XL U13393 ( .A(n5726), .B(n3757), .Z(n5792) );
  CNR2XL U13394 ( .A(n5722), .B(n3757), .Z(n5788) );
  CNR2X1 U13395 ( .A(n5171), .B(n3757), .Z(n5238) );
  CNR2X1 U13396 ( .A(n5745), .B(n3757), .Z(n5811) );
  CNR2X1 U13397 ( .A(n4722), .B(n3757), .Z(n4797) );
  CNR2X1 U13398 ( .A(n4746), .B(n3757), .Z(n4776) );
  CNR2X1 U13399 ( .A(n6169), .B(n3757), .Z(n6204) );
  CNR2X1 U13400 ( .A(n6153), .B(n3757), .Z(n6193) );
  CNR2X1 U13401 ( .A(n4534), .B(n3757), .Z(n6214) );
  CNR2X1 U13402 ( .A(n4570), .B(n3757), .Z(n6220) );
  CANR2X1 U13403 ( .A(mem_data1[486]), .B(n3898), .C(N8766), .D(n3681), .Z(
        n644) );
  CANR2X1 U13404 ( .A(mem_data1[480]), .B(n3898), .C(N8760), .D(n3680), .Z(
        n662) );
  CANR2X1 U13405 ( .A(mem_data1[481]), .B(n3898), .C(N8761), .D(n3680), .Z(
        n659) );
  CMXI2X1 U13406 ( .A0(n14057), .A1(n14030), .S(n3540), .Z(N8767) );
  CANR2X1 U13407 ( .A(mem_data1[352]), .B(n3898), .C(N8632), .D(n3680), .Z(
        n1046) );
  CMXI2X1 U13408 ( .A0(n13786), .A1(n13792), .S(n3750), .Z(n13799) );
  CANR2XL U13409 ( .A(N2324), .B(n3605), .C(n3638), .D(N8031), .Z(n1360) );
  CANR2X1 U13410 ( .A(mem_data1[238]), .B(n3898), .C(N8518), .D(n3679), .Z(
        n1388) );
  CMX2XL U13411 ( .A0(N8032), .A1(N8031), .S(n4243), .Z(n10112) );
  CANR2X1 U13412 ( .A(mem_data1[296]), .B(n3898), .C(N8576), .D(n3679), .Z(
        n1214) );
  CND2X1 U13413 ( .A(n5163), .B(n3213), .Z(n5230) );
  CMXI2X1 U13414 ( .A0(n13846), .A1(n13852), .S(n3750), .Z(n13858) );
  CANR2X1 U13415 ( .A(mem_data1[351]), .B(n3898), .C(N8631), .D(n3680), .Z(
        n1049) );
  CANR2X1 U13416 ( .A(mem_data1[484]), .B(n3898), .C(N8764), .D(n3680), .Z(
        n650) );
  CANR2X1 U13417 ( .A(mem_data1[483]), .B(n3898), .C(N8763), .D(n3680), .Z(
        n653) );
  CANR2X1 U13418 ( .A(mem_data1[485]), .B(n3898), .C(N8765), .D(n3680), .Z(
        n647) );
  CANR2X1 U13419 ( .A(mem_data1[369]), .B(n3898), .C(N8649), .D(n3680), .Z(
        n995) );
  CANR2X1 U13420 ( .A(N2564), .B(n3604), .C(n3638), .D(N7791), .Z(n640) );
  CMX2XL U13421 ( .A0(N7791), .A1(N7790), .S(n4280), .Z(n10921) );
  CEOX1 U13422 ( .A(N506), .B(mem_data1[488]), .Z(N7791) );
  CEOX1 U13423 ( .A(N266), .B(mem_data1[248]), .Z(N8031) );
  CND2X1 U13424 ( .A(n5172), .B(n3203), .Z(n5239) );
  CANR2X1 U13425 ( .A(mem_data1[356]), .B(n3898), .C(N8636), .D(n3680), .Z(
        n1034) );
  CANR2X1 U13426 ( .A(mem_data1[282]), .B(n3898), .C(n3678), .D(N8562), .Z(
        n1256) );
  CANR2X1 U13427 ( .A(mem_data1[298]), .B(n3898), .C(N8578), .D(n3679), .Z(
        n1208) );
  CANR2X1 U13428 ( .A(mem_data1[367]), .B(n3898), .C(N8647), .D(n3681), .Z(
        n1001) );
  CANR2X1 U13429 ( .A(N2436), .B(n3604), .C(n3637), .D(N7919), .Z(n1024) );
  CMX2XL U13430 ( .A0(N7919), .A1(N7918), .S(n4260), .Z(n10491) );
  CEOX1 U13431 ( .A(N378), .B(mem_data1[360]), .Z(N7919) );
  CMXI2X1 U13432 ( .A0(n13977), .A1(n13983), .S(n3750), .Z(n13990) );
  CANR2XL U13433 ( .A(N2448), .B(n3605), .C(n3638), .D(N7907), .Z(n988) );
  CMX2XL U13434 ( .A0(N7907), .A1(N7906), .S(n4260), .Z(n10533) );
  CEOX1 U13435 ( .A(N390), .B(mem_data1[372]), .Z(N7907) );
  CANR2X1 U13436 ( .A(mem_data1[286]), .B(n3898), .C(n3678), .D(N8566), .Z(
        n1244) );
  CANR2XL U13437 ( .A(N2571), .B(n3605), .C(n3638), .D(N7784), .Z(n619) );
  CMX2XL U13438 ( .A0(N7784), .A1(N7783), .S(n4236), .Z(n10945) );
  CEOX1 U13439 ( .A(N513), .B(mem_data1[495]), .Z(N7784) );
  CANR2X1 U13440 ( .A(N2327), .B(n3604), .C(n3638), .D(N8028), .Z(n1351) );
  CMX2XL U13441 ( .A0(N8029), .A1(N8028), .S(n4243), .Z(n10121) );
  CMXI2X1 U13442 ( .A0(n13352), .A1(n13346), .S(n4186), .Z(n3744) );
  CANR2X1 U13443 ( .A(mem_data1[300]), .B(n3898), .C(N8580), .D(n3679), .Z(
        n1202) );
  CANR2XL U13444 ( .A(N2568), .B(n3605), .C(n3638), .D(N7787), .Z(n628) );
  CMX2XL U13445 ( .A0(N7787), .A1(N7786), .S(n4231), .Z(n10936) );
  CND2X1 U13446 ( .A(n5213), .B(n3212), .Z(n5314) );
  CANR2X1 U13447 ( .A(mem_data1[355]), .B(n3898), .C(N8635), .D(n3681), .Z(
        n1037) );
  CMXI2X1 U13448 ( .A0(n13358), .A1(n13367), .S(n3750), .Z(n13374) );
  CANR2XL U13449 ( .A(N2467), .B(n3605), .C(n3638), .D(N7888), .Z(n931) );
  CANR2X1 U13450 ( .A(mem_data1[391]), .B(n3898), .C(N8671), .D(n3681), .Z(
        n929) );
  CMX2XL U13451 ( .A0(N7889), .A1(N7888), .S(n4258), .Z(n10590) );
  CMX2XL U13452 ( .A0(N7888), .A1(N7887), .S(n4258), .Z(n10593) );
  CANR2X1 U13453 ( .A(mem_data1[301]), .B(n3898), .C(N8581), .D(n3679), .Z(
        n1199) );
  CANR2X1 U13454 ( .A(mem_data1[429]), .B(n3898), .C(N8709), .D(n3682), .Z(
        n815) );
  CANR2XL U13455 ( .A(N2403), .B(n3604), .C(n3638), .D(N7952), .Z(n1123) );
  CANR2X1 U13456 ( .A(mem_data1[321]), .B(n3898), .C(N8601), .D(n3679), .Z(
        n1139) );
  CMX2XL U13457 ( .A0(N7953), .A1(N7952), .S(n4230), .Z(n10380) );
  CMX2XL U13458 ( .A0(N7952), .A1(N7951), .S(n4251), .Z(n10383) );
  CANR2X1 U13459 ( .A(mem_data1[428]), .B(n3898), .C(N8708), .D(n3679), .Z(
        n818) );
  CANR2XL U13460 ( .A(N2439), .B(n3605), .C(n3638), .D(N7916), .Z(n1015) );
  CMX2XL U13461 ( .A0(N7916), .A1(N7915), .S(n4256), .Z(n10503) );
  CEOX1 U13462 ( .A(N381), .B(mem_data1[363]), .Z(N7916) );
  CANR2XL U13463 ( .A(N2339), .B(n3605), .C(n3638), .D(N8016), .Z(n1315) );
  CANR2X1 U13464 ( .A(mem_data1[261]), .B(n3898), .C(N8541), .D(n3680), .Z(
        n1319) );
  CMX2XL U13465 ( .A0(N8017), .A1(N8016), .S(n4242), .Z(n10163) );
  CMX2XL U13466 ( .A0(N8016), .A1(N8015), .S(n4242), .Z(n10166) );
  CANR2XL U13467 ( .A(N2511), .B(n3605), .C(n3639), .D(N7844), .Z(n799) );
  CMX2XL U13468 ( .A0(N7845), .A1(N7844), .S(n4234), .Z(n10744) );
  CMX2XL U13469 ( .A0(N7844), .A1(N7843), .S(n4233), .Z(n10747) );
  CMXI2X1 U13470 ( .A0(n13361), .A1(n13370), .S(n3750), .Z(n13377) );
  CMXI2X1 U13471 ( .A0(n13798), .A1(n13804), .S(n3750), .Z(n13814) );
  CANR2X1 U13472 ( .A(mem_data1[426]), .B(n3898), .C(N8706), .D(n3682), .Z(
        n824) );
  CANR2X1 U13473 ( .A(mem_data1[427]), .B(n3898), .C(N8707), .D(n3682), .Z(
        n821) );
  CANR2X1 U13474 ( .A(mem_data1[376]), .B(n3898), .C(N8656), .D(n3681), .Z(
        n974) );
  CANR2XL U13475 ( .A(N2375), .B(n3605), .C(n3638), .D(N7980), .Z(n1207) );
  CANR2X1 U13476 ( .A(mem_data1[297]), .B(n3898), .C(N8577), .D(n3679), .Z(
        n1211) );
  CMX2XL U13477 ( .A0(N7981), .A1(N7980), .S(n4240), .Z(n10280) );
  CMX2XL U13478 ( .A0(N7980), .A1(N7979), .S(n4240), .Z(n10283) );
  CANR2X1 U13479 ( .A(mem_data1[425]), .B(n3898), .C(N8705), .D(n3682), .Z(
        n827) );
  CANR2X1 U13480 ( .A(mem_data1[249]), .B(n3898), .C(N8529), .D(n3680), .Z(
        n1355) );
  CEOX1 U13481 ( .A(N269), .B(mem_data1[251]), .Z(N8028) );
  CND2X1 U13482 ( .A(n5178), .B(n3203), .Z(n5245) );
  CANR2X1 U13483 ( .A(mem_data1[326]), .B(n3898), .C(N8606), .D(n3679), .Z(
        n1124) );
  CANR2X1 U13484 ( .A(mem_data1[388]), .B(n3898), .C(N8668), .D(n3681), .Z(
        n938) );
  CANR2X1 U13485 ( .A(mem_data1[324]), .B(n3898), .C(N8604), .D(n3679), .Z(
        n1130) );
  CANR2X1 U13486 ( .A(mem_data1[327]), .B(n3898), .C(N8607), .D(n3679), .Z(
        n1121) );
  CANR2XL U13487 ( .A(N2531), .B(n3605), .C(n3639), .D(N7824), .Z(n739) );
  CANR2X1 U13488 ( .A(mem_data1[455]), .B(n3898), .C(N8735), .D(n3680), .Z(
        n737) );
  CMX2XL U13489 ( .A0(N7825), .A1(N7824), .S(n4255), .Z(n10810) );
  CMX2XL U13490 ( .A0(N7824), .A1(N7823), .S(n4255), .Z(n10813) );
  CANR2X1 U13491 ( .A(mem_data1[386]), .B(n3898), .C(N8666), .D(n3681), .Z(
        n944) );
  CANR2X1 U13492 ( .A(mem_data1[389]), .B(n3898), .C(N8669), .D(n3681), .Z(
        n935) );
  CANR2X1 U13493 ( .A(mem_data1[325]), .B(n3898), .C(N8605), .D(n3679), .Z(
        n1127) );
  CANR2XL U13494 ( .A(N2337), .B(n3605), .C(n3638), .D(N8018), .Z(n1321) );
  CANR2X1 U13495 ( .A(mem_data1[259]), .B(n3898), .C(N8539), .D(n3680), .Z(
        n1325) );
  CMX2XL U13496 ( .A0(N8019), .A1(N8018), .S(n4242), .Z(n10154) );
  CMX2XL U13497 ( .A0(N8018), .A1(N8017), .S(n4242), .Z(n10157) );
  CANR2X1 U13498 ( .A(mem_data1[387]), .B(n3898), .C(N8667), .D(n3681), .Z(
        n941) );
  CANR2XL U13499 ( .A(N2509), .B(n3605), .C(n3639), .D(N7846), .Z(n805) );
  CMX2XL U13500 ( .A0(N7847), .A1(N7846), .S(n4236), .Z(n10738) );
  CMX2XL U13501 ( .A0(N7846), .A1(N7845), .S(n4235), .Z(n10741) );
  CANR2XL U13502 ( .A(N2366), .B(n3605), .C(n3638), .D(N7989), .Z(n1234) );
  CANR2X1 U13503 ( .A(mem_data1[279]), .B(n3898), .C(N8559), .D(n3679), .Z(
        n1265) );
  CMX2XL U13504 ( .A0(N7990), .A1(N7989), .S(n4244), .Z(n10250) );
  CMX2XL U13505 ( .A0(N7989), .A1(N7988), .S(n4245), .Z(n10253) );
  CANR2XL U13506 ( .A(N2443), .B(n3605), .C(n3638), .D(N7912), .Z(n1003) );
  CMX2XL U13507 ( .A0(N7912), .A1(N7911), .S(n4239), .Z(n10515) );
  CMX2XL U13508 ( .A0(N7913), .A1(N7912), .S(n4287), .Z(n10512) );
  CEOX1 U13509 ( .A(N385), .B(mem_data1[367]), .Z(N7912) );
  CMX2XL U13510 ( .A0(N7788), .A1(N7787), .S(n4280), .Z(n10930) );
  CMX2XL U13511 ( .A0(N7789), .A1(N7788), .S(n4230), .Z(n10927) );
  CEOX1 U13512 ( .A(N509), .B(mem_data1[491]), .Z(N7788) );
  CANR2X1 U13513 ( .A(mem_data1[430]), .B(n3898), .C(n3679), .D(N8710), .Z(
        n812) );
  CANR2XL U13514 ( .A(N2382), .B(n3605), .C(n3638), .D(N7973), .Z(n1186) );
  CANR2X1 U13515 ( .A(mem_data1[304]), .B(n3898), .C(N8584), .D(n3679), .Z(
        n1190) );
  CMX2XL U13516 ( .A0(N7974), .A1(N7973), .S(n4239), .Z(n10304) );
  CMX2XL U13517 ( .A0(N7973), .A1(N7972), .S(n4239), .Z(n10307) );
  CND2X1 U13518 ( .A(n5159), .B(n3201), .Z(n5226) );
  CANR2X1 U13519 ( .A(mem_data1[432]), .B(n3898), .C(N8712), .D(n3682), .Z(
        n806) );
  CANR2X1 U13520 ( .A(N2447), .B(n3604), .C(n3637), .D(N7908), .Z(n991) );
  CMX2XL U13521 ( .A0(N7908), .A1(N7907), .S(n4260), .Z(n10527) );
  CMX2XL U13522 ( .A0(N7909), .A1(N7908), .S(n4260), .Z(n10524) );
  CEOX1 U13523 ( .A(N389), .B(mem_data1[371]), .Z(N7908) );
  CANR2X1 U13524 ( .A(mem_data1[433]), .B(n3898), .C(n3678), .D(N8713), .Z(
        n803) );
  CMX2XL U13525 ( .A0(N8036), .A1(N8035), .S(n4244), .Z(n10100) );
  CMX2XL U13526 ( .A0(N8037), .A1(N8036), .S(n4244), .Z(n10097) );
  CEOX1 U13527 ( .A(N261), .B(mem_data1[243]), .Z(N8036) );
  CANR2X1 U13528 ( .A(mem_data1[431]), .B(n3898), .C(N8711), .D(n3682), .Z(
        n809) );
  CANR2XL U13529 ( .A(N2529), .B(n3605), .C(n3639), .D(N7826), .Z(n745) );
  CANR2X1 U13530 ( .A(mem_data1[450]), .B(n3898), .C(N8730), .D(n3680), .Z(
        n752) );
  CMX2XL U13531 ( .A0(N7827), .A1(N7826), .S(n4255), .Z(n10804) );
  CMX2XL U13532 ( .A0(N7826), .A1(N7825), .S(n4255), .Z(n10807) );
  CANR2X1 U13533 ( .A(mem_data1[453]), .B(n3898), .C(N8733), .D(n3679), .Z(
        n743) );
  CANR2XL U13534 ( .A(N2570), .B(n3605), .C(n3638), .D(N7785), .Z(n622) );
  CMX2XL U13535 ( .A0(N7786), .A1(N7785), .S(n4231), .Z(n10939) );
  CMX2XL U13536 ( .A0(N7785), .A1(N7784), .S(n4254), .Z(n10942) );
  CND2X1 U13537 ( .A(n5217), .B(n3214), .Z(n5318) );
  CANR2XL U13538 ( .A(N2321), .B(n3605), .C(n3638), .D(N8034), .Z(n1369) );
  CMX2XL U13539 ( .A0(N8035), .A1(N8034), .S(n4243), .Z(n10103) );
  CMX2XL U13540 ( .A0(N8034), .A1(N8033), .S(n4243), .Z(n10106) );
  CND2X1 U13541 ( .A(n5165), .B(n3207), .Z(n5232) );
  CANR2XL U13542 ( .A(N2401), .B(n3604), .C(n3638), .D(N7954), .Z(n1129) );
  CANR2X1 U13543 ( .A(mem_data1[323]), .B(n3898), .C(N8603), .D(n3679), .Z(
        n1133) );
  CMX2XL U13544 ( .A0(N7955), .A1(N7954), .S(n4250), .Z(n10374) );
  CMX2XL U13545 ( .A0(N7954), .A1(N7953), .S(n4236), .Z(n10377) );
  CANR2X1 U13546 ( .A(mem_data1[451]), .B(n3898), .C(N8731), .D(n3679), .Z(
        n749) );
  CANR2XL U13547 ( .A(N2441), .B(n3605), .C(n3638), .D(N7914), .Z(n1009) );
  CMX2XL U13548 ( .A0(N7915), .A1(N7914), .S(n4260), .Z(n10506) );
  CMX2XL U13549 ( .A0(N7914), .A1(N7913), .S(n4240), .Z(n10509) );
  CND2X1 U13550 ( .A(n5215), .B(n3210), .Z(n5316) );
  CANR2XL U13551 ( .A(N2438), .B(n3605), .C(n3638), .D(N7917), .Z(n1018) );
  CMX2XL U13552 ( .A0(N7918), .A1(N7917), .S(n4287), .Z(n10494) );
  CMX2XL U13553 ( .A0(N7917), .A1(N7916), .S(n4243), .Z(n10500) );
  CND2X1 U13554 ( .A(n5207), .B(n3208), .Z(n5310) );
  CANR2XL U13555 ( .A(N2445), .B(n3605), .C(n3638), .D(N7910), .Z(n997) );
  CMX2XL U13556 ( .A0(N7910), .A1(N7909), .S(n4260), .Z(n10521) );
  CMX2XL U13557 ( .A0(N7911), .A1(N7910), .S(n4240), .Z(n10518) );
  CEOX1 U13558 ( .A(N387), .B(mem_data1[369]), .Z(N7910) );
  CANR2XL U13559 ( .A(N2454), .B(n3605), .C(n3638), .D(N7901), .Z(n970) );
  CMX2XL U13560 ( .A0(N7902), .A1(N7901), .S(n4260), .Z(n10548) );
  CMX2XL U13561 ( .A0(N7901), .A1(N7900), .S(n4260), .Z(n10551) );
  CND2X1 U13562 ( .A(n5176), .B(n3211), .Z(n5243) );
  CND2X1 U13563 ( .A(n5169), .B(n3207), .Z(n5237) );
  CMXI2X1 U13564 ( .A0(n5087), .A1(n5030), .S(n4221), .Z(n5127) );
  CND2X1 U13565 ( .A(n5205), .B(n3208), .Z(n5308) );
  CANR2XL U13566 ( .A(N2317), .B(n3605), .C(n3638), .D(N8038), .Z(n1381) );
  CMX2XL U13567 ( .A0(N8038), .A1(N8037), .S(n4244), .Z(n10091) );
  CMX2XL U13568 ( .A0(N8039), .A1(N8038), .S(n4244), .Z(n10088) );
  CEOX1 U13569 ( .A(N259), .B(mem_data1[241]), .Z(N8038) );
  CANR2XL U13570 ( .A(N2494), .B(n3604), .C(n3638), .D(N7861), .Z(n850) );
  CANR2X1 U13571 ( .A(mem_data1[416]), .B(n3898), .C(N8696), .D(n3681), .Z(
        n854) );
  CMX2XL U13572 ( .A0(N7862), .A1(N7861), .S(n4256), .Z(n10687) );
  CMX2XL U13573 ( .A0(N7861), .A1(N7860), .S(n4256), .Z(n10690) );
  CANR2XL U13574 ( .A(N2325), .B(n3605), .C(n3638), .D(N8030), .Z(n1357) );
  CMX2XL U13575 ( .A0(N8031), .A1(N8030), .S(n4243), .Z(n10115) );
  CMX2XL U13576 ( .A0(N8030), .A1(N8029), .S(n4243), .Z(n10118) );
  CND2X1 U13577 ( .A(n5174), .B(n3207), .Z(n5241) );
  CNR2X1 U13578 ( .A(n3762), .B(n5081), .Z(n5150) );
  CND2X1 U13579 ( .A(n5199), .B(n3200), .Z(n5301) );
  CND2X1 U13580 ( .A(n3712), .B(n3205), .Z(n5235) );
  CND2X1 U13581 ( .A(n5150), .B(n3201), .Z(n5218) );
  CANR2XL U13582 ( .A(N2489), .B(n3605), .C(n3638), .D(n3714), .Z(n865) );
  CMX2XL U13583 ( .A0(n3714), .A1(N7865), .S(n4256), .Z(n10675) );
  CMX2XL U13584 ( .A0(N7867), .A1(n3714), .S(n4256), .Z(n10672) );
  CMXI2X1 U13585 ( .A0(n4968), .A1(n4994), .S(n3896), .Z(n5023) );
  CANR2X1 U13586 ( .A(mem_data1[412]), .B(n3898), .C(N8692), .D(n3681), .Z(
        n866) );
  CMXI2XL U13587 ( .A0(n4732), .A1(n4731), .S(n3763), .Z(n3745) );
  CMXI2X1 U13588 ( .A0(n4659), .A1(n4660), .S(n3752), .Z(n4731) );
  CANR2X1 U13589 ( .A(mem_data1[410]), .B(n3898), .C(N8690), .D(n3681), .Z(
        n872) );
  CANR2XL U13590 ( .A(N2523), .B(n3605), .C(n3639), .D(N7832), .Z(n763) );
  CMX2XL U13591 ( .A0(N7833), .A1(N7832), .S(n4279), .Z(n10783) );
  CMX2XL U13592 ( .A0(N7832), .A1(N7831), .S(n4280), .Z(n10786) );
  CMXI2XL U13593 ( .A0(n13788), .A1(n13815), .S(n3532), .Z(N8693) );
  CANR2XL U13594 ( .A(N2361), .B(n3605), .C(n3638), .D(N7994), .Z(n1249) );
  CANR2X1 U13595 ( .A(mem_data1[283]), .B(n3898), .C(N8563), .D(n3680), .Z(
        n1253) );
  CMX2XL U13596 ( .A0(N7995), .A1(N7994), .S(n4239), .Z(n10235) );
  CMX2XL U13597 ( .A0(N7994), .A1(N7993), .S(n4245), .Z(n10238) );
  CANR2X1 U13598 ( .A(mem_data1[411]), .B(n3898), .C(N8691), .D(n3681), .Z(
        n869) );
  CANR2XL U13599 ( .A(N2331), .B(n3605), .C(n3638), .D(N8024), .Z(n1339) );
  CMX2XL U13600 ( .A0(N8024), .A1(N8023), .S(n4242), .Z(n10139) );
  CANR2XL U13601 ( .A(N2558), .B(n3605), .C(n3639), .D(N7797), .Z(n658) );
  CMX2XL U13602 ( .A0(N7797), .A1(N7796), .S(n4232), .Z(n10903) );
  CMX2XL U13603 ( .A0(N7798), .A1(N7797), .S(n4228), .Z(n10897) );
  CEOX1 U13604 ( .A(N500), .B(mem_data1[482]), .Z(N7797) );
  CND2X1 U13605 ( .A(n5482), .B(n4394), .Z(n4560) );
  CND2X1 U13606 ( .A(N5601), .B(n3698), .Z(n774) );
  CANR2X1 U13607 ( .A(mem_data1[112]), .B(n3898), .C(n3678), .D(N8392), .Z(
        n1766) );
  CANR2X1 U13608 ( .A(mem_data1[110]), .B(n3898), .C(N8390), .D(n3679), .Z(
        n1772) );
  CANR2X1 U13609 ( .A(mem_data1[118]), .B(n3898), .C(N8398), .D(n3680), .Z(
        n1748) );
  CANR2XL U13610 ( .A(N2553), .B(n3605), .C(n3639), .D(N7802), .Z(n673) );
  CANR2X1 U13611 ( .A(mem_data1[477]), .B(n3898), .C(N8757), .D(n3680), .Z(
        n671) );
  CMX2XL U13612 ( .A0(N7803), .A1(N7802), .S(n4253), .Z(n10882) );
  CMX2XL U13613 ( .A0(N7802), .A1(N7801), .S(n4253), .Z(n10885) );
  CANR2XL U13614 ( .A(N2308), .B(n3605), .C(n3638), .D(N8047), .Z(n1408) );
  CMX2XL U13615 ( .A0(N8047), .A1(N8046), .S(n4245), .Z(n10064) );
  CEOX1 U13616 ( .A(N250), .B(mem_data1[232]), .Z(N8047) );
  CANR2XL U13617 ( .A(N2425), .B(n3604), .C(n3638), .D(N7930), .Z(n1057) );
  CANR2X1 U13618 ( .A(mem_data1[347]), .B(n3898), .C(N8627), .D(n3680), .Z(
        n1061) );
  CMX2XL U13619 ( .A0(N7931), .A1(N7930), .S(n4237), .Z(n10452) );
  CMX2XL U13620 ( .A0(N7930), .A1(N7929), .S(n4237), .Z(n10455) );
  CANR2X1 U13621 ( .A(mem_data1[475]), .B(n3898), .C(N8755), .D(n3680), .Z(
        n677) );
  CMXI2X1 U13622 ( .A0(n12741), .A1(n12749), .S(n3750), .Z(n12755) );
  CANR2XL U13623 ( .A(N2395), .B(n3604), .C(n3638), .D(N7960), .Z(n1147) );
  CMX2XL U13624 ( .A0(N7961), .A1(N7960), .S(n4252), .Z(n10353) );
  CMX2XL U13625 ( .A0(N7960), .A1(N7959), .S(n4235), .Z(n10356) );
  CMXI2X1 U13626 ( .A0(n13418), .A1(n13384), .S(n3540), .Z(N8575) );
  CANR2XL U13627 ( .A(N2499), .B(n3604), .C(n3638), .D(N7856), .Z(n835) );
  CANR2X1 U13628 ( .A(mem_data1[423]), .B(n3898), .C(N8703), .D(n3682), .Z(
        n833) );
  CMX2XL U13629 ( .A0(N7856), .A1(N7855), .S(n4279), .Z(n10708) );
  CANR2XL U13630 ( .A(N2369), .B(n3605), .C(n3638), .D(N7986), .Z(n1225) );
  CMXI2X1 U13631 ( .A0(n12807), .A1(n12783), .S(n3541), .Z(N8397) );
  CANR2XL U13632 ( .A(N2459), .B(n3605), .C(n3638), .D(N7896), .Z(n955) );
  CMX2XL U13633 ( .A0(N7896), .A1(N7895), .S(n4259), .Z(n10569) );
  CMX2XL U13634 ( .A0(N7897), .A1(N7896), .S(n4259), .Z(n10566) );
  CMXI2X1 U13635 ( .A0(n13337), .A1(n13343), .S(n3750), .Z(n13350) );
  CANR2X1 U13636 ( .A(mem_data1[421]), .B(n3898), .C(N8701), .D(n3682), .Z(
        n839) );
  CANR2XL U13637 ( .A(N2137), .B(n3605), .C(n3638), .D(N8218), .Z(n1921) );
  CMX2XL U13638 ( .A0(N8218), .A1(N8217), .S(n4255), .Z(n10999) );
  CANR2XL U13639 ( .A(N2434), .B(n3604), .C(n3638), .D(N7921), .Z(n1030) );
  CEOX1 U13640 ( .A(N376), .B(mem_data1[358]), .Z(N7921) );
  CANR2XL U13641 ( .A(N2265), .B(n3605), .C(n3639), .D(N8090), .Z(n1537) );
  CANR2X1 U13642 ( .A(mem_data1[181]), .B(n3898), .C(N8461), .D(n3681), .Z(
        n1559) );
  CMX2XL U13643 ( .A0(N8091), .A1(N8090), .S(n4249), .Z(n9911) );
  CMX2XL U13644 ( .A0(N8090), .A1(N8089), .S(n4249), .Z(n9914) );
  CANR2X1 U13645 ( .A(mem_data1[182]), .B(n3898), .C(N8462), .D(n3681), .Z(
        n1556) );
  CANR2X1 U13646 ( .A(mem_data1[59]), .B(n3898), .C(N8339), .D(n3679), .Z(
        n1925) );
  CANR2X1 U13647 ( .A(mem_data1[228]), .B(n3898), .C(N8508), .D(n3679), .Z(
        n1418) );
  CEOX1 U13648 ( .A(N248), .B(mem_data1[230]), .Z(N8049) );
  CND2X1 U13649 ( .A(N5452), .B(n3698), .Z(n1221) );
  CMXI2X1 U13650 ( .A0(n12745), .A1(n12751), .S(n3750), .Z(n12761) );
  CMXI2X1 U13651 ( .A0(n4558), .A1(n4559), .S(N2066), .Z(n4600) );
  CANR2X1 U13652 ( .A(mem_data1[183]), .B(n3898), .C(N8463), .D(n3681), .Z(
        n1553) );
  CMXI2X1 U13653 ( .A0(n12725), .A1(n12726), .S(n3750), .Z(n12743) );
  CMXI2X1 U13654 ( .A0(n12786), .A1(n12762), .S(n3541), .Z(N8390) );
  CANR2X1 U13655 ( .A(mem_data1[111]), .B(n3898), .C(N8391), .D(n3680), .Z(
        n1769) );
  CANR2X1 U13656 ( .A(mem_data1[113]), .B(n3898), .C(N8393), .D(n3680), .Z(
        n1763) );
  CANR2XL U13657 ( .A(N2562), .B(n3605), .C(n3638), .D(N7793), .Z(n646) );
  CMX2XL U13658 ( .A0(N7793), .A1(N7792), .S(n4280), .Z(n10915) );
  CEOX1 U13659 ( .A(N504), .B(mem_data1[486]), .Z(N7793) );
  CMXI2X1 U13660 ( .A0(n12732), .A1(n12733), .S(n3750), .Z(n12747) );
  CANR2XL U13661 ( .A(N2498), .B(n3604), .C(n3638), .D(N7857), .Z(n838) );
  CMX2XL U13662 ( .A0(N7857), .A1(N7856), .S(n4255), .Z(n10705) );
  CANR2XL U13663 ( .A(N2370), .B(n3604), .C(n3638), .D(N7985), .Z(n1222) );
  CANR2X1 U13664 ( .A(mem_data1[294]), .B(n3898), .C(N8574), .D(n3679), .Z(
        n1220) );
  CMX2XL U13665 ( .A0(N7986), .A1(N7985), .S(n4239), .Z(n10265) );
  CMX2XL U13666 ( .A0(N7985), .A1(N7984), .S(n4240), .Z(n10268) );
  CANR2X1 U13667 ( .A(mem_data1[187]), .B(n3898), .C(N8467), .D(n3681), .Z(
        n1541) );
  CIVXL U13668 ( .A(n4646), .Z(n3746) );
  CND2X1 U13669 ( .A(n5040), .B(n4398), .Z(n5049) );
  CND2XL U13670 ( .A(n5048), .B(n4399), .Z(n5056) );
  CANR2XL U13671 ( .A(N2563), .B(n3605), .C(n3638), .D(N7792), .Z(n643) );
  CMX2XL U13672 ( .A0(N7792), .A1(N7791), .S(n4228), .Z(n10918) );
  CANR2XL U13673 ( .A(N2368), .B(n3605), .C(n3638), .D(N7987), .Z(n1228) );
  CMX2XL U13674 ( .A0(N7988), .A1(N7987), .S(n4243), .Z(n10256) );
  CMX2XL U13675 ( .A0(N7987), .A1(N7986), .S(n4240), .Z(n10262) );
  CND2X1 U13676 ( .A(n5195), .B(n3212), .Z(n5297) );
  CNR2X1 U13677 ( .A(n5162), .B(n3758), .Z(n5229) );
  CANR2X1 U13678 ( .A(mem_data1[291]), .B(n3898), .C(N8571), .D(n3679), .Z(
        n1229) );
  CANR2XL U13679 ( .A(N2497), .B(n3604), .C(n3638), .D(N7858), .Z(n841) );
  CANR2X1 U13680 ( .A(mem_data1[419]), .B(n3898), .C(N8699), .D(n3681), .Z(
        n845) );
  CMX2XL U13681 ( .A0(N7859), .A1(N7858), .S(n4249), .Z(n10696) );
  CMX2XL U13682 ( .A0(N7858), .A1(N7857), .S(n4249), .Z(n10699) );
  CANR2XL U13683 ( .A(N2435), .B(n3604), .C(n3638), .D(N7920), .Z(n1027) );
  CMX2XL U13684 ( .A0(N7921), .A1(N7920), .S(n4261), .Z(n10485) );
  CMX2XL U13685 ( .A0(N7920), .A1(N7919), .S(n4243), .Z(n10488) );
  CMXI2XL U13686 ( .A0(n3219), .A1(n4643), .S(n3764), .Z(n3748) );
  CMXI2XL U13687 ( .A0(n4643), .A1(n4646), .S(n4221), .Z(n4690) );
  CANR2XL U13688 ( .A(N2329), .B(n3605), .C(n3638), .D(N8026), .Z(n1345) );
  CMXI2X1 U13689 ( .A0(n4724), .A1(n4723), .S(n3763), .Z(n3749) );
  CND2X1 U13690 ( .A(n5193), .B(n3214), .Z(n5295) );
  CNR2X1 U13691 ( .A(n5160), .B(n3757), .Z(n5227) );
  CANR2XL U13692 ( .A(N2561), .B(n3605), .C(n3639), .D(N7794), .Z(n649) );
  CMX2XL U13693 ( .A0(N7795), .A1(N7794), .S(n4229), .Z(n10909) );
  CMX2XL U13694 ( .A0(N7794), .A1(N7793), .S(n4233), .Z(n10912) );
  CMXI2X1 U13695 ( .A0(n4515), .A1(n4516), .S(n3896), .Z(n4646) );
  CANR2XL U13696 ( .A(N2433), .B(n3605), .C(n3638), .D(N7922), .Z(n1033) );
  CMX2XL U13697 ( .A0(N7923), .A1(N7922), .S(n4261), .Z(n10479) );
  CMX2XL U13698 ( .A0(N7922), .A1(N7921), .S(n4261), .Z(n10482) );
  CANR2XL U13699 ( .A(N2430), .B(n3605), .C(n3638), .D(N7925), .Z(n1042) );
  CMX2XL U13700 ( .A0(N7926), .A1(N7925), .S(n4237), .Z(n10470) );
  CMX2XL U13701 ( .A0(N7925), .A1(N7924), .S(n4239), .Z(n10473) );
  CND2X1 U13702 ( .A(n5191), .B(n3210), .Z(n5293) );
  CANR2X1 U13703 ( .A(mem_data1[185]), .B(n3898), .C(N8465), .D(n3681), .Z(
        n1547) );
  CANR2XL U13704 ( .A(N2136), .B(n3605), .C(n3638), .D(N8219), .Z(n1924) );
  CMX2XL U13705 ( .A0(N8220), .A1(N8219), .S(n4253), .Z(n10933) );
  CMX2XL U13706 ( .A0(N8219), .A1(N8218), .S(n4230), .Z(n10966) );
  CANR2XL U13707 ( .A(N2393), .B(n3604), .C(n3638), .D(N7962), .Z(n1153) );
  CMX2XL U13708 ( .A0(N7963), .A1(N7962), .S(n4279), .Z(n10347) );
  CMX2XL U13709 ( .A0(N7962), .A1(N7961), .S(n4253), .Z(n10350) );
  CANR2XL U13710 ( .A(N2521), .B(n3605), .C(n3639), .D(N7834), .Z(n769) );
  CMX2XL U13711 ( .A0(N7835), .A1(N7834), .S(n4235), .Z(n10777) );
  CMX2XL U13712 ( .A0(N7834), .A1(N7833), .S(n4228), .Z(n10780) );
  CANR2XL U13713 ( .A(N2457), .B(n3605), .C(n3638), .D(N7898), .Z(n961) );
  CMX2XL U13714 ( .A0(N7899), .A1(N7898), .S(n4259), .Z(n10557) );
  CMX2XL U13715 ( .A0(N7898), .A1(N7897), .S(n4259), .Z(n10560) );
  CND2X1 U13716 ( .A(n4959), .B(n4397), .Z(n4966) );
  CND2X1 U13717 ( .A(n6250), .B(n3740), .Z(n6352) );
  CNR2IX1 U13718 ( .B(n6183), .A(n3215), .Z(n6250) );
  CANR2XL U13719 ( .A(N2328), .B(n3605), .C(n3638), .D(N8027), .Z(n1348) );
  CMX2XL U13720 ( .A0(N8028), .A1(N8027), .S(n4243), .Z(n10124) );
  CMX2XL U13721 ( .A0(N8027), .A1(N8026), .S(n4243), .Z(n10130) );
  CANR2XL U13722 ( .A(N2330), .B(n3605), .C(n3638), .D(N8025), .Z(n1342) );
  CMX2XL U13723 ( .A0(N8026), .A1(N8025), .S(n4243), .Z(n10133) );
  CMX2XL U13724 ( .A0(N8025), .A1(N8024), .S(n4242), .Z(n10136) );
  CND2X1 U13725 ( .A(n5184), .B(n3209), .Z(n5251) );
  CMXI2XL U13726 ( .A0(n4600), .A1(n4603), .S(n3194), .Z(n4619) );
  CND2X1 U13727 ( .A(n5497), .B(n4394), .Z(n4559) );
  CMXI2X1 U13728 ( .A0(n12769), .A1(n12775), .S(lenin0[1]), .Z(n12782) );
  CANR2X1 U13729 ( .A(mem_data1[120]), .B(n3898), .C(N8400), .D(n3680), .Z(
        n1742) );
  CEOX1 U13730 ( .A(N140), .B(mem_data1[122]), .Z(N8157) );
  CNR2X1 U13731 ( .A(n3763), .B(n4715), .Z(n4655) );
  CANR2XL U13732 ( .A(N2179), .B(n3605), .C(n3638), .D(N8176), .Z(n1795) );
  CEOX1 U13733 ( .A(N121), .B(mem_data1[103]), .Z(N8176) );
  CMXI2X1 U13734 ( .A0(n13058), .A1(n13034), .S(n3542), .Z(N8470) );
  CANR2X1 U13735 ( .A(mem_data1[189]), .B(n3898), .C(N8469), .D(n3681), .Z(
        n1535) );
  CMXI2X1 U13736 ( .A0(n13061), .A1(n13037), .S(n3542), .Z(N8471) );
  CANR2XL U13737 ( .A(N2139), .B(n3605), .C(n3638), .D(N8216), .Z(n1915) );
  CANR2X1 U13738 ( .A(mem_data1[61]), .B(n3898), .C(N8341), .D(n3679), .Z(
        n1919) );
  CMX2XL U13739 ( .A0(N8217), .A1(N8216), .S(n4252), .Z(n11036) );
  CMX2XL U13740 ( .A0(N8216), .A1(N8215), .S(n4251), .Z(n11069) );
  CND2XL U13741 ( .A(n6056), .B(n4412), .Z(n6061) );
  CMXI2X1 U13742 ( .A0(n12986), .A1(n12992), .S(n3750), .Z(n13003) );
  CEOX1 U13743 ( .A(N138), .B(mem_data1[120]), .Z(N8159) );
  CND2X1 U13744 ( .A(n4610), .B(n3892), .Z(n4707) );
  CNR2X1 U13745 ( .A(n4219), .B(n4517), .Z(n4645) );
  CANR2XL U13746 ( .A(N2191), .B(n3605), .C(n3639), .D(N8164), .Z(n1759) );
  CMX2XL U13747 ( .A0(N8165), .A1(N8164), .S(n4286), .Z(n9655) );
  CMX2XL U13748 ( .A0(N8164), .A1(N8163), .S(n4286), .Z(n9662) );
  CEOX1 U13749 ( .A(N133), .B(mem_data1[115]), .Z(N8164) );
  CANR2XL U13750 ( .A(N2307), .B(n3605), .C(n3638), .D(N8048), .Z(n1411) );
  CMX2XL U13751 ( .A0(N8049), .A1(N8048), .S(n4245), .Z(n10055) );
  CMX2XL U13752 ( .A0(N8048), .A1(N8047), .S(n4245), .Z(n10058) );
  CANR2XL U13753 ( .A(N2197), .B(n3605), .C(n3638), .D(N8158), .Z(n1741) );
  CMX2XL U13754 ( .A0(N8159), .A1(N8158), .S(n4285), .Z(n9679) );
  CMX2XL U13755 ( .A0(N8158), .A1(N8157), .S(n4285), .Z(n9682) );
  CNR2X1 U13756 ( .A(n3764), .B(n3700), .Z(n4761) );
  CANR2XL U13757 ( .A(N2178), .B(n3605), .C(n3639), .D(N8177), .Z(n1798) );
  CMX2XL U13758 ( .A0(N8178), .A1(N8177), .S(n4286), .Z(n12271) );
  CMX2XL U13759 ( .A0(N8177), .A1(N8176), .S(n4287), .Z(n9649) );
  CNR2XL U13760 ( .A(n4696), .B(n3758), .Z(n4785) );
  CND2X1 U13761 ( .A(n5553), .B(n4392), .Z(n4548) );
  CND2X1 U13762 ( .A(n5576), .B(n4392), .Z(n4547) );
  CND2X1 U13763 ( .A(n5560), .B(n4392), .Z(n4549) );
  CND2X1 U13764 ( .A(n5569), .B(n4392), .Z(n4546) );
  CND2X1 U13765 ( .A(n5583), .B(n4392), .Z(n4544) );
  CND2X1 U13766 ( .A(n5590), .B(n4392), .Z(n4545) );
  CND2X1 U13767 ( .A(n5597), .B(n4392), .Z(n4542) );
  CANR2XL U13768 ( .A(N2199), .B(n3605), .C(n3638), .D(N8156), .Z(n1735) );
  CMX2XL U13769 ( .A0(N8157), .A1(N8156), .S(n4285), .Z(n9688) );
  CMX2XL U13770 ( .A0(N8156), .A1(N8155), .S(n4285), .Z(n9691) );
  CNR2X1 U13771 ( .A(n3764), .B(n3706), .Z(n4705) );
  CMXI2XL U13772 ( .A0(n4601), .A1(n4600), .S(n3188), .Z(n4639) );
  CMXI2XL U13773 ( .A0(n4598), .A1(n4601), .S(n3190), .Z(n4616) );
  CANR2XL U13774 ( .A(N2201), .B(n3605), .C(n3638), .D(N8154), .Z(n1729) );
  CANR2X1 U13775 ( .A(mem_data1[115]), .B(n3898), .C(N8395), .D(n3680), .Z(
        n1757) );
  CMX2XL U13776 ( .A0(N8155), .A1(N8154), .S(n4285), .Z(n9694) );
  CND2X1 U13777 ( .A(n5528), .B(n4393), .Z(n4552) );
  CND2X1 U13778 ( .A(n5546), .B(n4393), .Z(n4551) );
  CND2X1 U13779 ( .A(n5534), .B(n4393), .Z(n4553) );
  CND2X1 U13780 ( .A(n5540), .B(n4393), .Z(n4550) );
  CND2X1 U13781 ( .A(n5510), .B(n4393), .Z(n4557) );
  CND2X1 U13782 ( .A(n5516), .B(n4393), .Z(n4554) );
  CND2X1 U13783 ( .A(n5522), .B(n4393), .Z(n4555) );
  CANR2X1 U13784 ( .A(mem_data1[405]), .B(n3898), .C(N8685), .D(n3681), .Z(
        n887) );
  CND2X1 U13785 ( .A(n5186), .B(n3215), .Z(n5253) );
  CNR2X1 U13786 ( .A(n3765), .B(n5088), .Z(n5153) );
  CND2X1 U13787 ( .A(n4975), .B(n3894), .Z(n5031) );
  CMXI2XL U13788 ( .A0(n5030), .A1(n4975), .S(n4222), .Z(n5088) );
  CND2X1 U13789 ( .A(n6056), .B(n4396), .Z(n4936) );
  CND2X1 U13790 ( .A(n4935), .B(n4396), .Z(n4942) );
  CND2X1 U13791 ( .A(n4941), .B(n4396), .Z(n4948) );
  CND2X1 U13792 ( .A(n6037), .B(n4396), .Z(n4918) );
  CND2X1 U13793 ( .A(n6041), .B(n4396), .Z(n4923) );
  CND2X1 U13794 ( .A(n6046), .B(n4396), .Z(n4927) );
  CND2X1 U13795 ( .A(n6051), .B(n4396), .Z(n4931) );
  CANR2X1 U13796 ( .A(mem_data1[123]), .B(n3898), .C(N8403), .D(n3680), .Z(
        n1733) );
  CEOX1 U13797 ( .A(N143), .B(mem_data1[125]), .Z(N8154) );
  CNR2X1 U13798 ( .A(n3766), .B(n4727), .Z(n4765) );
  CND2X1 U13799 ( .A(n4651), .B(n3894), .Z(n4693) );
  CMXI2XL U13800 ( .A0(n4652), .A1(n4651), .S(n4227), .Z(n4727) );
  CANR2XL U13801 ( .A(N2203), .B(n3605), .C(n3638), .D(N8152), .Z(n1723) );
  CMX2XL U13802 ( .A0(N8152), .A1(N8151), .S(n4284), .Z(n9703) );
  CND2X1 U13803 ( .A(n4665), .B(n3895), .Z(n4701) );
  CND2X1 U13804 ( .A(n5188), .B(n3206), .Z(n5291) );
  CNR2X1 U13805 ( .A(n5156), .B(n3759), .Z(n5223) );
  CNR2X1 U13806 ( .A(n5117), .B(n3896), .Z(n5144) );
  CND2X1 U13807 ( .A(n5055), .B(n4399), .Z(n5063) );
  CND2XL U13808 ( .A(n5062), .B(n4399), .Z(n5070) );
  CND2XL U13809 ( .A(n5069), .B(n4399), .Z(n5077) );
  CND2XL U13810 ( .A(n5090), .B(n4399), .Z(n5096) );
  CND2XL U13811 ( .A(n5076), .B(n4399), .Z(n5084) );
  CND2XL U13812 ( .A(n5083), .B(n4399), .Z(n5091) );
  CNR2X1 U13813 ( .A(n4741), .B(n3759), .Z(n4774) );
  CND2X1 U13814 ( .A(n4672), .B(n4224), .Z(n4710) );
  CND2X1 U13815 ( .A(n5611), .B(n4391), .Z(n4540) );
  CND2X1 U13816 ( .A(n5618), .B(n4391), .Z(n4541) );
  CND2X1 U13817 ( .A(n5625), .B(n4391), .Z(n4538) );
  CND2X1 U13818 ( .A(n5632), .B(n4391), .Z(n4539) );
  CND2X1 U13819 ( .A(n5654), .B(n4391), .Z(n4535) );
  CND2X1 U13820 ( .A(n5640), .B(n4391), .Z(n4536) );
  CND2X1 U13821 ( .A(n5647), .B(n4391), .Z(n4537) );
  CIVXL U13822 ( .A(wr_ptr[9]), .Z(n4414) );
  CIVXL U13823 ( .A(wr_ptr[9]), .Z(n4401) );
  CIVXL U13824 ( .A(wr_ptr[9]), .Z(n4402) );
  CIVXL U13825 ( .A(wr_ptr[9]), .Z(n4403) );
  CND2X1 U13826 ( .A(n6252), .B(n3739), .Z(n6354) );
  CIVX1 U13827 ( .A(n4390), .Z(n4388) );
  CND2X1 U13828 ( .A(n6248), .B(n3736), .Z(n6350) );
  CNR2X1 U13829 ( .A(n3828), .B(n6023), .Z(N751) );
  CNR2X1 U13830 ( .A(n3822), .B(n5920), .Z(N658) );
  CNR2X1 U13831 ( .A(n3826), .B(n6348), .Z(N1020) );
  CNR2X1 U13832 ( .A(n3833), .B(n6492), .Z(N1001) );
  CNR2X1 U13833 ( .A(n3820), .B(n6458), .Z(N972) );
  CNR2X1 U13834 ( .A(n3821), .B(n5991), .Z(N722) );
  CNR2X1 U13835 ( .A(n3823), .B(n6022), .Z(N750) );
  CNR2X1 U13836 ( .A(n3839), .B(n5856), .Z(N78) );
  CIVXL U13837 ( .A(n13401), .Z(n4432) );
  CANR2XL U13838 ( .A(N2180), .B(n3605), .C(n3639), .D(N8175), .Z(n1792) );
  CANR2X1 U13839 ( .A(mem_data1[94]), .B(n3898), .C(N8374), .D(n3680), .Z(
        n1820) );
  CMX2XL U13840 ( .A0(N8176), .A1(N8175), .S(n4286), .Z(n9656) );
  CMX2XL U13841 ( .A0(N8175), .A1(N8174), .S(n4288), .Z(n9650) );
  CANR2X1 U13842 ( .A(mem_data1[102]), .B(n3898), .C(N8382), .D(n3680), .Z(
        n1796) );
  CEOX1 U13843 ( .A(N122), .B(mem_data1[104]), .Z(N8175) );
  CND2X1 U13844 ( .A(n4607), .B(n4224), .Z(n4706) );
  CNR2X1 U13845 ( .A(n4510), .B(n3896), .Z(n4642) );
  CNR2X1 U13846 ( .A(n3242), .B(n3758), .Z(n4780) );
  CANR2XL U13847 ( .A(N2202), .B(n3605), .C(n3638), .D(N8153), .Z(n1726) );
  CMX2XL U13848 ( .A0(N8154), .A1(N8153), .S(n4284), .Z(n9697) );
  CMX2XL U13849 ( .A0(N8153), .A1(N8152), .S(n4284), .Z(n9700) );
  CNR2X1 U13850 ( .A(n3763), .B(n4731), .Z(n4769) );
  CND2XL U13851 ( .A(n4991), .B(n4395), .Z(n4999) );
  CND2X1 U13852 ( .A(n6032), .B(n4395), .Z(n4915) );
  CND2X1 U13853 ( .A(n5469), .B(n4395), .Z(n4565) );
  CND2X1 U13854 ( .A(n6029), .B(n4395), .Z(n4912) );
  CND2X1 U13855 ( .A(n5466), .B(n4395), .Z(n4564) );
  CND2X1 U13856 ( .A(n6027), .B(n4395), .Z(n4910) );
  CND2X1 U13857 ( .A(n5464), .B(n4395), .Z(n4566) );
  CAN3X1 U13858 ( .A(wr_ptr[6]), .B(n3199), .C(wr_ptr[7]), .Z(n3751) );
  CIVX1 U13859 ( .A(n4414), .Z(n4400) );
  CANR2X1 U13860 ( .A(mem_data1[162]), .B(n3898), .C(N8442), .D(n3681), .Z(
        n1616) );
  CNR2X1 U13861 ( .A(n3834), .B(n5326), .Z(N54) );
  CNR2X1 U13862 ( .A(n3819), .B(n5326), .Z(N182) );
  CANR2XL U13863 ( .A(N6223), .B(n3605), .C(n3193), .D(n3639), .Z(n2122) );
  CANR2XL U13864 ( .A(N6223), .B(n2105), .C(n3191), .D(n3898), .Z(n2123) );
  CANR2X1 U13865 ( .A(mem_data1[186]), .B(n3898), .C(N8466), .D(n3681), .Z(
        n1544) );
  CNR2X1 U13866 ( .A(n3765), .B(n4723), .Z(n4743) );
  CND2XL U13867 ( .A(n5475), .B(n3193), .Z(n5485) );
  CND2XL U13868 ( .A(n5471), .B(n3189), .Z(n5480) );
  CND2XL U13869 ( .A(n4916), .B(n3195), .Z(n4925) );
  CND2XL U13870 ( .A(n4913), .B(n3195), .Z(n4920) );
  CND2XL U13871 ( .A(n4587), .B(n3189), .Z(n4630) );
  CND2XL U13872 ( .A(n4604), .B(n3191), .Z(n4620) );
  CND2XL U13873 ( .A(n6039), .B(n3191), .Z(n6049) );
  CND2XL U13874 ( .A(n6034), .B(n3193), .Z(n6044) );
  CFA1XL U13875 ( .A(n3189), .B(lenin0[1]), .CI(\r347/carry [1]), .CO(
        \r347/carry [2]), .S(N6223) );
  CNIVXL U13876 ( .A(N2069), .Z(n3752) );
  CNIVX1 U13877 ( .A(n4436), .Z(n4211) );
  CNR2X1 U13878 ( .A(n3845), .B(n5503), .Z(N66) );
  CNR2X1 U13879 ( .A(n3824), .B(n5503), .Z(N194) );
  CIVDX1 U13880 ( .A(N2070), .Z0(n3755), .Z1(n3756) );
  CNIVX1 U13881 ( .A(n3755), .Z(n3763) );
  CNIVX1 U13882 ( .A(n3755), .Z(n3764) );
  CNIVX1 U13883 ( .A(n3755), .Z(n3765) );
  CNIVX1 U13884 ( .A(n3755), .Z(n3766) );
  CIVXL U13885 ( .A(n4376), .Z(n3767) );
  CIVXL U13886 ( .A(n4376), .Z(n3768) );
  CNIVX3 U13887 ( .A(n3770), .Z(n3771) );
  CNIVX2 U13888 ( .A(n3770), .Z(n3772) );
  CNIVX2 U13889 ( .A(n3770), .Z(n3773) );
  CNIVX2 U13890 ( .A(n4305), .Z(n3774) );
  CNIVX2 U13891 ( .A(n3767), .Z(n3775) );
  CNIVX2 U13892 ( .A(n3767), .Z(n3776) );
  CNIVX2 U13893 ( .A(n4306), .Z(n3777) );
  CNIVX1 U13894 ( .A(n3769), .Z(n3778) );
  CNIVX1 U13895 ( .A(n3769), .Z(n3779) );
  CNIVX1 U13896 ( .A(n3769), .Z(n3780) );
  CNIVX1 U13897 ( .A(n3769), .Z(n3781) );
  CNIVX1 U13898 ( .A(n3780), .Z(n3782) );
  CNIVX1 U13899 ( .A(n3778), .Z(n3783) );
  CNIVX1 U13900 ( .A(n3779), .Z(n3784) );
  CNIVX1 U13901 ( .A(n3781), .Z(n3785) );
  CIVDX1 U13902 ( .A(n3767), .Z0(n3786), .Z1(n3787) );
  CIVDX1 U13903 ( .A(n3767), .Z0(n3788), .Z1(n3789) );
  CNIVX2 U13904 ( .A(n3787), .Z(n3790) );
  CNIVX2 U13905 ( .A(n3787), .Z(n3791) );
  CNIVX2 U13906 ( .A(n3787), .Z(n3792) );
  CNIVX2 U13907 ( .A(n3787), .Z(n3793) );
  CNIVX2 U13908 ( .A(n3789), .Z(n3794) );
  CNIVX2 U13909 ( .A(n3789), .Z(n3795) );
  CNIVX2 U13910 ( .A(n3789), .Z(n3796) );
  CNIVX2 U13911 ( .A(n3789), .Z(n3797) );
  CNIVX1 U13912 ( .A(n3786), .Z(n3798) );
  CNIVX1 U13913 ( .A(n3786), .Z(n3799) );
  CNIVX1 U13914 ( .A(n3786), .Z(n3800) );
  CNIVX1 U13915 ( .A(n3786), .Z(n3801) );
  CIVDX1 U13916 ( .A(n3768), .Z0(n3802), .Z1(n3803) );
  CIVDX1 U13917 ( .A(n3768), .Z0(n3218), .Z1(n3804) );
  CNIVX2 U13918 ( .A(n3803), .Z(n3805) );
  CNIVX2 U13919 ( .A(n3803), .Z(n3806) );
  CNIVX2 U13920 ( .A(n3803), .Z(n3807) );
  CNIVX2 U13921 ( .A(n3803), .Z(n3808) );
  CNIVX2 U13922 ( .A(n3804), .Z(n3809) );
  CNIVX2 U13923 ( .A(n3804), .Z(n3810) );
  CNIVX2 U13924 ( .A(n3804), .Z(n3811) );
  CNIVX2 U13925 ( .A(n3804), .Z(n3812) );
  CNIVX1 U13926 ( .A(n4385), .Z(n4376) );
  CNIVX1 U13927 ( .A(n4385), .Z(n4377) );
  CNIVX1 U13928 ( .A(n4385), .Z(n4378) );
  CANR2XL U13929 ( .A(N6227), .B(n2105), .C(n3898), .D(n3213), .Z(n2115) );
  CNR2IXL U13930 ( .B(n6185), .A(n3203), .Z(n6252) );
  CNR2IXL U13931 ( .B(n6180), .A(n3211), .Z(n6248) );
  CNIVX1 U13932 ( .A(n3814), .Z(n3815) );
  CNIVX1 U13933 ( .A(n3814), .Z(n3816) );
  CNIVX1 U13934 ( .A(n3814), .Z(n3817) );
  CNIVX1 U13935 ( .A(n3814), .Z(n3818) );
  CNIVX1 U13936 ( .A(n3814), .Z(n3819) );
  CNIVX1 U13937 ( .A(n3814), .Z(n3820) );
  CNIVX1 U13938 ( .A(n3814), .Z(n3821) );
  CNIVX1 U13939 ( .A(n3814), .Z(n3822) );
  CNIVX1 U13940 ( .A(n3814), .Z(n3823) );
  CNIVX1 U13941 ( .A(n3814), .Z(n3824) );
  CNIVX1 U13942 ( .A(n3814), .Z(n3825) );
  CNIVX1 U13943 ( .A(n3814), .Z(n3826) );
  CNIVX1 U13944 ( .A(n3814), .Z(n3827) );
  CNIVX1 U13945 ( .A(n3814), .Z(n3828) );
  CNIVX1 U13946 ( .A(n3814), .Z(n3829) );
  CNIVX1 U13947 ( .A(n3814), .Z(n3830) );
  CNIVX1 U13948 ( .A(n3814), .Z(n3831) );
  CNIVX1 U13949 ( .A(n3814), .Z(n3832) );
  CNIVX1 U13950 ( .A(n3814), .Z(n3833) );
  CNIVX1 U13951 ( .A(n3813), .Z(n3834) );
  CNIVX1 U13952 ( .A(n3813), .Z(n3835) );
  CNIVX1 U13953 ( .A(n3813), .Z(n3836) );
  CNIVX1 U13954 ( .A(n3813), .Z(n3837) );
  CNIVX1 U13955 ( .A(n3813), .Z(n3838) );
  CNIVX1 U13956 ( .A(n3813), .Z(n3839) );
  CNIVX1 U13957 ( .A(n3813), .Z(n3840) );
  CNIVX1 U13958 ( .A(n3813), .Z(n3841) );
  CNIVX1 U13959 ( .A(n3813), .Z(n3842) );
  CNIVX1 U13960 ( .A(n3813), .Z(n3843) );
  CNIVX1 U13961 ( .A(n3813), .Z(n3844) );
  CNIVX1 U13962 ( .A(n3813), .Z(n3845) );
  CNIVX1 U13963 ( .A(n3813), .Z(n3846) );
  CNIVX1 U13964 ( .A(n3813), .Z(n3847) );
  CNIVX1 U13965 ( .A(n3813), .Z(n3848) );
  CNIVX1 U13966 ( .A(n3813), .Z(n3849) );
  CNIVX1 U13967 ( .A(n3813), .Z(n3850) );
  CNIVX1 U13968 ( .A(n3813), .Z(n3851) );
  CNIVX1 U13969 ( .A(n3813), .Z(n3852) );
  CNIVX1 U13970 ( .A(n3813), .Z(n3853) );
  CIVDXL U13971 ( .A(lenin0[0]), .Z0(n3854), .Z1(n3855) );
  CIVDXL U13972 ( .A(lenin0[0]), .Z0(n3856), .Z1(n3857) );
  CIVDXL U13973 ( .A(lenin0[0]), .Z0(n3858), .Z1(n3859) );
  CIVDXL U13974 ( .A(lenin0[0]), .Z0(n3860), .Z1(n3861) );
  CNIVX3 U13975 ( .A(n3855), .Z(n3862) );
  CNIVX3 U13976 ( .A(n3855), .Z(n3863) );
  CNIVX3 U13977 ( .A(n3855), .Z(n3864) );
  CNIVX3 U13978 ( .A(n3855), .Z(n3865) );
  CNIVX3 U13979 ( .A(n3855), .Z(n3866) );
  CNIVX3 U13980 ( .A(n3857), .Z(n3867) );
  CNIVX3 U13981 ( .A(n3857), .Z(n3868) );
  CNIVX3 U13982 ( .A(n3857), .Z(n3869) );
  CNIVX3 U13983 ( .A(n3857), .Z(n3870) );
  CNIVX3 U13984 ( .A(n3857), .Z(n3871) );
  CNIVX3 U13985 ( .A(n3859), .Z(n3872) );
  CNIVX3 U13986 ( .A(n3859), .Z(n3873) );
  CNIVX3 U13987 ( .A(n3859), .Z(n3874) );
  CNIVX3 U13988 ( .A(n3859), .Z(n3875) );
  CNIVX3 U13989 ( .A(n3859), .Z(n3876) );
  CNIVX3 U13990 ( .A(n3861), .Z(n3877) );
  CNIVX3 U13991 ( .A(n3861), .Z(n3878) );
  CNIVX3 U13992 ( .A(n3861), .Z(n3879) );
  CNIVX3 U13993 ( .A(n3861), .Z(n3880) );
  CNIVX3 U13994 ( .A(n3861), .Z(n3881) );
  CNIVX1 U13995 ( .A(n3854), .Z(n3882) );
  CNIVX1 U13996 ( .A(n3854), .Z(n3883) );
  CNIVX1 U13997 ( .A(n3854), .Z(n3884) );
  CNIVX1 U13998 ( .A(n3854), .Z(n3885) );
  CNIVX1 U13999 ( .A(n3854), .Z(n3886) );
  CNIVX1 U14000 ( .A(n3856), .Z(n3887) );
  CNIVX1 U14001 ( .A(n3856), .Z(n3888) );
  CNIVX1 U14002 ( .A(n3858), .Z(n3889) );
  CNIVX1 U14003 ( .A(n3860), .Z(n3890) );
  CNIVX1 U14004 ( .A(n4302), .Z(n4301) );
  CIVX2 U14005 ( .A(n4390), .Z(n4389) );
  CIVXL U14006 ( .A(n3754), .Z(n4221) );
  CIVXL U14007 ( .A(n3754), .Z(n4222) );
  CIVXL U14008 ( .A(n3754), .Z(n4223) );
  CIVXL U14009 ( .A(n3754), .Z(n4224) );
  CIVXL U14010 ( .A(n3754), .Z(n4225) );
  CIVXL U14011 ( .A(n4301), .Z(n4294) );
  CIVX1 U14012 ( .A(lenin0[0]), .Z(n4302) );
  CIVX1 U14013 ( .A(lenin0[0]), .Z(n4303) );
  CIVX1 U14014 ( .A(lenin0[0]), .Z(n4304) );
  CIVX2 U14015 ( .A(lenin0[2]), .Z(n4385) );
  CIVXL U14016 ( .A(n4390), .Z(n4386) );
  CIVXL U14017 ( .A(n4390), .Z(n4387) );
  CIVXL U14018 ( .A(n4413), .Z(n4391) );
  CIVXL U14019 ( .A(n4413), .Z(n4392) );
  CIVXL U14020 ( .A(n4405), .Z(n4393) );
  CIVXL U14021 ( .A(n4405), .Z(n4394) );
  CIVXL U14022 ( .A(n4405), .Z(n4395) );
  CIVXL U14023 ( .A(n4404), .Z(n4396) );
  CIVXL U14024 ( .A(n4404), .Z(n4397) );
  CIVXL U14025 ( .A(n4409), .Z(n4398) );
  CIVXL U14026 ( .A(n4409), .Z(n4399) );
  CIVX2 U14027 ( .A(wr_ptr[9]), .Z(n4404) );
  CIVX2 U14028 ( .A(wr_ptr[9]), .Z(n4405) );
  CIVX2 U14029 ( .A(wr_ptr[9]), .Z(n4406) );
  CIVX2 U14030 ( .A(wr_ptr[9]), .Z(n4407) );
  CIVX2 U14031 ( .A(wr_ptr[9]), .Z(n4408) );
  CIVX2 U14032 ( .A(wr_ptr[9]), .Z(n4409) );
  CIVX2 U14033 ( .A(wr_ptr[9]), .Z(n4410) );
  CIVX2 U14034 ( .A(wr_ptr[9]), .Z(n4411) );
  CIVX2 U14035 ( .A(wr_ptr[9]), .Z(n4412) );
  CIVX2 U14036 ( .A(wr_ptr[9]), .Z(n4413) );
  CENX1 U14037 ( .A(N3108), .B(\r349/carry [8]), .Z(N6230) );
  COR2X1 U14038 ( .A(N3106), .B(N3105), .Z(\r349/carry [7]) );
  CENX1 U14039 ( .A(N3106), .B(N3105), .Z(N6228) );
  CENX1 U14040 ( .A(n4400), .B(\sub_84/carry [9]), .Z(N2075) );
  COR2X1 U14041 ( .A(n4386), .B(\sub_84/carry [8]), .Z(\sub_84/carry [9]) );
  CENX1 U14042 ( .A(n4389), .B(\sub_84/carry [8]), .Z(N2074) );
  COR2X1 U14043 ( .A(n3816), .B(\sub_84/carry [7]), .Z(\sub_84/carry [8]) );
  CENX1 U14044 ( .A(n3817), .B(\sub_84/carry [7]), .Z(N2073) );
  COR2X1 U14045 ( .A(n3724), .B(n3209), .Z(\sub_84/carry [7]) );
  CENX1 U14046 ( .A(n3725), .B(n3211), .Z(N2072) );
  CEOX1 U14047 ( .A(n4389), .B(\r347/carry [8]), .Z(N3108) );
  CAN2X1 U14048 ( .A(\r347/carry [7]), .B(n3815), .Z(\r347/carry [8]) );
  CAN2X1 U14049 ( .A(\r347/carry [6]), .B(n3723), .Z(\r347/carry [7]) );
  CEOX1 U14050 ( .A(n3722), .B(\r347/carry [6]), .Z(N3106) );
  CAN2X1 U14051 ( .A(\r347/carry [5]), .B(n3205), .Z(\r347/carry [6]) );
  CEOX1 U14052 ( .A(n3207), .B(\r347/carry [5]), .Z(N3105) );
  CEOX1 U14053 ( .A(n3758), .B(\r347/carry [4]), .Z(N6226) );
  CEOX1 U14054 ( .A(n3870), .B(N2066), .Z(N6222) );
  CIVX2 U14055 ( .A(N3105), .Z(N6227) );
  CIVX2 U14056 ( .A(n7930), .Z(n4416) );
  CIVX2 U14057 ( .A(n8598), .Z(n4417) );
  CIVX2 U14058 ( .A(n8932), .Z(n4418) );
  CIVX2 U14059 ( .A(n8264), .Z(n4419) );
  CIVX2 U14060 ( .A(n11002), .Z(n4420) );
  CIVX2 U14061 ( .A(n11670), .Z(n4421) );
  CIVX2 U14062 ( .A(n12004), .Z(n4422) );
  CIVX2 U14063 ( .A(n11336), .Z(n4423) );
  CIVX2 U14064 ( .A(n14741), .Z(n4425) );
  CIVX2 U14065 ( .A(n7257), .Z(n4429) );
  CIVX2 U14066 ( .A(n7594), .Z(n4430) );
  CIVX2 U14067 ( .A(n10666), .Z(n4431) );
  CIVX2 U14068 ( .A(n13738), .Z(n4433) );
  CIVX2 U14069 ( .A(pushin0), .Z(n4434) );
  CIVX2 U14070 ( .A(reqin0), .Z(n4435) );
  CIVX2 U14071 ( .A(lenout[3]), .Z(n4438) );
  CIVX2 U14072 ( .A(lenout[2]), .Z(n4439) );
  CMXI2X1 U14073 ( .A0(n4535), .A1(n4537), .S(n4210), .Z(n4572) );
  CMXI2X1 U14074 ( .A0(n4536), .A1(n4539), .S(n4206), .Z(n4574) );
  CMXI2X1 U14075 ( .A0(n4572), .A1(n4574), .S(n3188), .Z(n4510) );
  CMXI2X1 U14076 ( .A0(n4538), .A1(n4541), .S(n4204), .Z(n4573) );
  CMXI2X1 U14077 ( .A0(n4540), .A1(n4543), .S(n4203), .Z(n4576) );
  CMXI2X1 U14078 ( .A0(n4573), .A1(n4576), .S(n3190), .Z(n4512) );
  CMXI2X1 U14079 ( .A0(n4510), .A1(n4512), .S(n4218), .Z(n4607) );
  CMXI2X1 U14080 ( .A0(n4542), .A1(n4545), .S(n4203), .Z(n4575) );
  CMXI2X1 U14081 ( .A0(n4544), .A1(n4547), .S(n4204), .Z(n4578) );
  CMXI2X1 U14082 ( .A0(n4575), .A1(n4578), .S(n3192), .Z(n4511) );
  CMXI2X1 U14083 ( .A0(n4546), .A1(n4549), .S(n4208), .Z(n4577) );
  CMXI2X1 U14084 ( .A0(n4548), .A1(n4551), .S(n4209), .Z(n4580) );
  CMXI2X1 U14085 ( .A0(n4577), .A1(n4580), .S(n3190), .Z(n4514) );
  CMXI2X1 U14086 ( .A0(n4511), .A1(n4514), .S(n4217), .Z(n4609) );
  CMXI2X1 U14087 ( .A0(n4607), .A1(n4609), .S(n4227), .Z(n4668) );
  CMXI2X1 U14088 ( .A0(n4550), .A1(n4553), .S(n4210), .Z(n4579) );
  CMXI2X1 U14089 ( .A0(n4552), .A1(n4555), .S(n4204), .Z(n4582) );
  CMXI2X1 U14090 ( .A0(n4579), .A1(n4582), .S(n3190), .Z(n4513) );
  CMXI2X1 U14091 ( .A0(n4554), .A1(n4557), .S(n4205), .Z(n4581) );
  CMXI2X1 U14092 ( .A0(n4556), .A1(n4559), .S(n4208), .Z(n4584) );
  CMXI2X1 U14093 ( .A0(n4581), .A1(n4584), .S(n3194), .Z(n4516) );
  CMXI2X1 U14094 ( .A0(n4513), .A1(n4516), .S(n4218), .Z(n4608) );
  CMXI2X1 U14095 ( .A0(n4558), .A1(n4561), .S(n4203), .Z(n4583) );
  CMXI2X1 U14096 ( .A0(n4560), .A1(n4563), .S(n4204), .Z(n4586) );
  CMXI2X1 U14097 ( .A0(n4562), .A1(n4565), .S(n4205), .Z(n4585) );
  CMXI2X1 U14098 ( .A0(n4564), .A1(n4566), .S(n4211), .Z(n4587) );
  CMXI2X1 U14099 ( .A0(n4585), .A1(n4587), .S(n3192), .Z(n4517) );
  CMXI2X1 U14100 ( .A0(n3710), .A1(n4517), .S(n4220), .Z(n4610) );
  CMXI2X1 U14101 ( .A0(n4608), .A1(n4610), .S(n4221), .Z(n4669) );
  CMXI2X1 U14102 ( .A0(n4668), .A1(n4669), .S(n3764), .Z(n4806) );
  CMXI2X1 U14103 ( .A0(n4441), .A1(n4443), .S(n4207), .Z(n4464) );
  CMXI2X1 U14104 ( .A0(n4442), .A1(n4445), .S(n4209), .Z(n4466) );
  CMXI2X1 U14105 ( .A0(n4464), .A1(n4466), .S(n3192), .Z(n4486) );
  CMXI2X1 U14106 ( .A0(n4444), .A1(n4447), .S(n4207), .Z(n4465) );
  CMXI2X1 U14107 ( .A0(n4446), .A1(n4449), .S(n4211), .Z(n4468) );
  CMXI2X1 U14108 ( .A0(n4465), .A1(n4468), .S(n3188), .Z(n4488) );
  CMXI2X1 U14109 ( .A0(n4486), .A1(n4488), .S(n4219), .Z(n4507) );
  CMXI2X1 U14110 ( .A0(n4448), .A1(n4451), .S(n4204), .Z(n4467) );
  CMXI2X1 U14111 ( .A0(n4450), .A1(n4453), .S(n4207), .Z(n4470) );
  CMXI2X1 U14112 ( .A0(n4467), .A1(n4470), .S(n3190), .Z(n4487) );
  CMXI2X1 U14113 ( .A0(n4452), .A1(n4455), .S(n4206), .Z(n4469) );
  CMXI2X1 U14114 ( .A0(n4454), .A1(n4457), .S(n4203), .Z(n4472) );
  CMXI2X1 U14115 ( .A0(n4469), .A1(n4472), .S(n3190), .Z(n4490) );
  CMXI2X1 U14116 ( .A0(n4487), .A1(n4490), .S(n4218), .Z(n4506) );
  CMXI2X1 U14117 ( .A0(n4456), .A1(n4459), .S(n4209), .Z(n4471) );
  CMXI2X1 U14118 ( .A0(n4458), .A1(n4461), .S(n4205), .Z(n4474) );
  CMXI2X1 U14119 ( .A0(n4471), .A1(n4474), .S(n3188), .Z(n4489) );
  CMXI2X1 U14120 ( .A0(n4460), .A1(n4463), .S(n4211), .Z(n4473) );
  CMXI2X1 U14121 ( .A0(n4462), .A1(n6062), .S(n4205), .Z(n6068) );
  CMXI2X1 U14122 ( .A0(n4473), .A1(n6068), .S(n3190), .Z(n6078) );
  CMXI2X1 U14123 ( .A0(n4489), .A1(n6078), .S(n4219), .Z(n6095) );
  CMXI2X1 U14124 ( .A0(n4506), .A1(n6095), .S(n4227), .Z(n6127) );
  CMXI2X1 U14125 ( .A0(n4531), .A1(n6127), .S(n3766), .Z(n6174) );
  CMXI2X1 U14126 ( .A0(n4443), .A1(n4442), .S(n4207), .Z(n4477) );
  CMXI2X1 U14127 ( .A0(n4475), .A1(n4477), .S(n3188), .Z(n4491) );
  CMXI2X1 U14128 ( .A0(n4445), .A1(n4444), .S(n4209), .Z(n4476) );
  CMXI2X1 U14129 ( .A0(n4447), .A1(n4446), .S(n4211), .Z(n4479) );
  CMXI2X1 U14130 ( .A0(n4476), .A1(n4479), .S(n3188), .Z(n4493) );
  CMXI2X1 U14131 ( .A0(n4491), .A1(n4493), .S(n4215), .Z(n4509) );
  CMXI2X1 U14132 ( .A0(n4449), .A1(n4448), .S(n4207), .Z(n4478) );
  CMXI2X1 U14133 ( .A0(n4451), .A1(n4450), .S(n4210), .Z(n4481) );
  CMXI2X1 U14134 ( .A0(n4478), .A1(n4481), .S(n3194), .Z(n4492) );
  CMXI2X1 U14135 ( .A0(n4453), .A1(n4452), .S(n4208), .Z(n4480) );
  CMXI2X1 U14136 ( .A0(n4455), .A1(n4454), .S(n4203), .Z(n4483) );
  CMXI2X1 U14137 ( .A0(n4480), .A1(n4483), .S(n3192), .Z(n4495) );
  CMXI2X1 U14138 ( .A0(n4492), .A1(n4495), .S(n4212), .Z(n4508) );
  CMXI2X1 U14139 ( .A0(n4457), .A1(n4456), .S(n4204), .Z(n4482) );
  CMXI2X1 U14140 ( .A0(n4459), .A1(n4458), .S(n4205), .Z(n4485) );
  CMXI2X1 U14141 ( .A0(n4482), .A1(n4485), .S(n3188), .Z(n4494) );
  CMXI2X1 U14142 ( .A0(n4461), .A1(n4460), .S(n4206), .Z(n4484) );
  CMXI2X1 U14143 ( .A0(n4463), .A1(n4462), .S(n4204), .Z(n6073) );
  CMXI2X1 U14144 ( .A0(n4484), .A1(n6073), .S(n3194), .Z(n6082) );
  CMXI2X1 U14145 ( .A0(n4494), .A1(n6082), .S(n4219), .Z(n6098) );
  CMXI2X1 U14146 ( .A0(n4508), .A1(n6098), .S(n4226), .Z(n6130) );
  CMXI2X1 U14147 ( .A0(n4532), .A1(n6130), .S(n3765), .Z(n6176) );
  CMXI2X1 U14148 ( .A0(n4466), .A1(n4465), .S(n3194), .Z(n4498) );
  CMXI2X1 U14149 ( .A0(n4496), .A1(n4498), .S(n3247), .Z(n4520) );
  CMXI2X1 U14150 ( .A0(n4468), .A1(n4467), .S(n3194), .Z(n4497) );
  CMXI2X1 U14151 ( .A0(n4470), .A1(n4469), .S(n3194), .Z(n4500) );
  CMXI2X1 U14152 ( .A0(n4497), .A1(n4500), .S(n4213), .Z(n4519) );
  CMXI2X1 U14153 ( .A0(n4472), .A1(n4471), .S(n3190), .Z(n4499) );
  CMXI2X1 U14154 ( .A0(n4474), .A1(n4473), .S(n3194), .Z(n6087) );
  CMXI2X1 U14155 ( .A0(n4499), .A1(n6087), .S(n4216), .Z(n6102) );
  CMXI2X1 U14156 ( .A0(n4519), .A1(n6102), .S(n4224), .Z(n6133) );
  CMXI2X1 U14157 ( .A0(n4477), .A1(n4476), .S(n3188), .Z(n4503) );
  CMXI2X1 U14158 ( .A0(n4501), .A1(n4503), .S(n4220), .Z(n4522) );
  CMXI2X1 U14159 ( .A0(n4479), .A1(n4478), .S(n3192), .Z(n4502) );
  CMXI2X1 U14160 ( .A0(n4481), .A1(n4480), .S(n3192), .Z(n4505) );
  CMXI2X1 U14161 ( .A0(n4502), .A1(n4505), .S(n4217), .Z(n4521) );
  CMXI2X1 U14162 ( .A0(n4483), .A1(n4482), .S(n3190), .Z(n4504) );
  CMXI2X1 U14163 ( .A0(n4485), .A1(n4484), .S(n3190), .Z(n6091) );
  CMXI2X1 U14164 ( .A0(n4504), .A1(n6091), .S(n4214), .Z(n6106) );
  CMXI2X1 U14165 ( .A0(n4521), .A1(n6106), .S(n4227), .Z(n6136) );
  CMXI2X1 U14166 ( .A0(n4534), .A1(n6136), .S(n3762), .Z(n6180) );
  CMXI2X1 U14167 ( .A0(n4488), .A1(n4487), .S(n3246), .Z(n4523) );
  CMXI2X1 U14168 ( .A0(n4490), .A1(n4489), .S(n4215), .Z(n6110) );
  CMXI2X1 U14169 ( .A0(n4523), .A1(n6110), .S(n4226), .Z(n6139) );
  CMXI2X1 U14170 ( .A0(n4568), .A1(n6139), .S(n3763), .Z(n6183) );
  CMXI2X1 U14171 ( .A0(n4493), .A1(n4492), .S(n4217), .Z(n4525) );
  CMXI2X1 U14172 ( .A0(n4495), .A1(n4494), .S(n4212), .Z(n6114) );
  CMXI2X1 U14173 ( .A0(n4525), .A1(n6114), .S(n4227), .Z(n6142) );
  CMXI2X1 U14174 ( .A0(n4569), .A1(n6142), .S(n3765), .Z(n6185) );
  CMXI2X1 U14175 ( .A0(n4498), .A1(n4497), .S(n3247), .Z(n4527) );
  CMXI2X1 U14176 ( .A0(n4500), .A1(n4499), .S(n4217), .Z(n6118) );
  CMXI2X1 U14177 ( .A0(n4527), .A1(n6118), .S(n4226), .Z(n6145) );
  CMXI2X1 U14178 ( .A0(n4570), .A1(n6145), .S(n3762), .Z(n6187) );
  CMXI2X1 U14179 ( .A0(n4503), .A1(n4502), .S(n4217), .Z(n4529) );
  CMXI2X1 U14180 ( .A0(n4505), .A1(n4504), .S(n4212), .Z(n6122) );
  CMXI2X1 U14181 ( .A0(n4529), .A1(n6122), .S(n4221), .Z(n6148) );
  CMXI2X1 U14182 ( .A0(n4571), .A1(n6148), .S(n3763), .Z(n6189) );
  CMXI2X1 U14183 ( .A0(n4507), .A1(n4506), .S(n4223), .Z(n6151) );
  CMXI2X1 U14184 ( .A0(n4509), .A1(n4508), .S(n4225), .Z(n6153) );
  CMXI2X1 U14185 ( .A0(n4512), .A1(n4511), .S(n4215), .Z(n4644) );
  CMXI2X1 U14186 ( .A0(n4514), .A1(n4513), .S(n4215), .Z(n4643) );
  CMXI2X1 U14187 ( .A0(n3746), .A1(n3748), .S(n3747), .Z(n4750) );
  CMXI2X1 U14188 ( .A0(n4917), .A1(n4518), .S(n3835), .Z(N118) );
  CMXI2X1 U14189 ( .A0(n4520), .A1(n4519), .S(n4226), .Z(n6157) );
  CMXI2X1 U14190 ( .A0(n4522), .A1(n4521), .S(n4226), .Z(n6160) );
  CMXI2X1 U14191 ( .A0(n4524), .A1(n4523), .S(n4226), .Z(n6163) );
  CMXI2X1 U14192 ( .A0(n4526), .A1(n4525), .S(n4225), .Z(n6166) );
  CMXI2X1 U14193 ( .A0(n4528), .A1(n4527), .S(n4226), .Z(n6169) );
  CMXI2X1 U14194 ( .A0(n4530), .A1(n4529), .S(n4224), .Z(n6172) );
  CMXI2X1 U14195 ( .A0(n4537), .A1(n4536), .S(n4208), .Z(n4591) );
  CMXI2X1 U14196 ( .A0(n4589), .A1(n4591), .S(n3192), .Z(n4613) );
  CMXI2X1 U14197 ( .A0(n4539), .A1(n4538), .S(n4210), .Z(n4590) );
  CMXI2X1 U14198 ( .A0(n4541), .A1(n4540), .S(n4208), .Z(n4593) );
  CMXI2X1 U14199 ( .A0(n4590), .A1(n4593), .S(n3188), .Z(n4612) );
  CMXI2X1 U14200 ( .A0(n4543), .A1(n4542), .S(n4210), .Z(n4592) );
  CMXI2X1 U14201 ( .A0(n4545), .A1(n4544), .S(n4209), .Z(n4595) );
  CMXI2X1 U14202 ( .A0(n4592), .A1(n4595), .S(n3190), .Z(n4615) );
  CMXI2X1 U14203 ( .A0(n4612), .A1(n4615), .S(n3246), .Z(n4650) );
  CMXI2X1 U14204 ( .A0(n4648), .A1(n4650), .S(n4226), .Z(n4692) );
  CMXI2X1 U14205 ( .A0(n4547), .A1(n4546), .S(n4206), .Z(n4594) );
  CMXI2X1 U14206 ( .A0(n4549), .A1(n4548), .S(n4207), .Z(n4597) );
  CMXI2X1 U14207 ( .A0(n4594), .A1(n4597), .S(n3192), .Z(n4614) );
  CMXI2X1 U14208 ( .A0(n4551), .A1(n4550), .S(n4211), .Z(n4596) );
  CMXI2X1 U14209 ( .A0(n4553), .A1(n4552), .S(n4205), .Z(n4599) );
  CMXI2X1 U14210 ( .A0(n4596), .A1(n4599), .S(n3192), .Z(n4617) );
  CMXI2X1 U14211 ( .A0(n4614), .A1(n4617), .S(n3247), .Z(n4649) );
  CMXI2X1 U14212 ( .A0(n4555), .A1(n4554), .S(n4205), .Z(n4598) );
  CMXI2X1 U14213 ( .A0(n4557), .A1(n4556), .S(n4203), .Z(n4601) );
  CMXI2X1 U14214 ( .A0(n4561), .A1(n4560), .S(n4204), .Z(n4603) );
  CMXI2X1 U14215 ( .A0(n4616), .A1(n4619), .S(n4220), .Z(n4652) );
  CMXI2X1 U14216 ( .A0(n4649), .A1(n4652), .S(n4223), .Z(n4694) );
  CMXI2X1 U14217 ( .A0(n4692), .A1(n4694), .S(n3766), .Z(n4752) );
  CMXI2X1 U14218 ( .A0(n4563), .A1(n4562), .S(n4206), .Z(n4602) );
  CMXI2X1 U14219 ( .A0(n4565), .A1(n4564), .S(n4203), .Z(n4605) );
  CMXI2X1 U14220 ( .A0(n4602), .A1(n4605), .S(n3192), .Z(n4618) );
  CMXI2X1 U14221 ( .A0(n4618), .A1(n4620), .S(n4218), .Z(n4651) );
  CMXI2X1 U14222 ( .A0(n4921), .A1(n4567), .S(n3836), .Z(N119) );
  CMXI2X1 U14223 ( .A0(n4574), .A1(n4573), .S(n3190), .Z(n4622) );
  CMXI2X1 U14224 ( .A0(n4576), .A1(n4575), .S(n3194), .Z(n4625) );
  CMXI2X1 U14225 ( .A0(n4578), .A1(n4577), .S(n3192), .Z(n4624) );
  CMXI2X1 U14226 ( .A0(n4580), .A1(n4579), .S(n3192), .Z(n4627) );
  CMXI2X1 U14227 ( .A0(n4582), .A1(n4581), .S(n3190), .Z(n4626) );
  CMXI2X1 U14228 ( .A0(n4584), .A1(n4583), .S(n3192), .Z(n4629) );
  CMXI2X1 U14229 ( .A0(n4626), .A1(n4629), .S(n4220), .Z(n4660) );
  CMXI2X1 U14230 ( .A0(n4657), .A1(n4660), .S(n4226), .Z(n4698) );
  CMXI2X1 U14231 ( .A0(n4696), .A1(n4698), .S(n3762), .Z(n4754) );
  CMXI2X1 U14232 ( .A0(n4586), .A1(n4585), .S(n3194), .Z(n4628) );
  CMXI2X1 U14233 ( .A0(n4628), .A1(n4630), .S(n4217), .Z(n4659) );
  CMXI2X1 U14234 ( .A0(n4926), .A1(n4588), .S(n3845), .Z(N120) );
  CMXI2X1 U14235 ( .A0(n4591), .A1(n4590), .S(n3188), .Z(n4632) );
  CMXI2X1 U14236 ( .A0(n4593), .A1(n4592), .S(n3190), .Z(n4635) );
  CMXI2X1 U14237 ( .A0(n4632), .A1(n4635), .S(n4217), .Z(n4664) );
  CMXI2X1 U14238 ( .A0(n4662), .A1(n4664), .S(n4225), .Z(n4700) );
  CMXI2X1 U14239 ( .A0(n4595), .A1(n4594), .S(n3194), .Z(n4634) );
  CMXI2X1 U14240 ( .A0(n4597), .A1(n4596), .S(n3188), .Z(n4637) );
  CMXI2X1 U14241 ( .A0(n4634), .A1(n4637), .S(n3247), .Z(n4663) );
  CMXI2X1 U14242 ( .A0(n4599), .A1(n4598), .S(n3192), .Z(n4636) );
  CMXI2X1 U14243 ( .A0(n4636), .A1(n4639), .S(n4213), .Z(n4666) );
  CMXI2X1 U14244 ( .A0(n4700), .A1(n4702), .S(n3764), .Z(n4756) );
  CMXI2X1 U14245 ( .A0(n4605), .A1(n4604), .S(n3190), .Z(n4640) );
  CMXI2X1 U14246 ( .A0(n4638), .A1(n4640), .S(n4218), .Z(n4665) );
  CMXI2X1 U14247 ( .A0(n4930), .A1(n4606), .S(n3846), .Z(N121) );
  CMXI2X1 U14248 ( .A0(n4609), .A1(n4608), .S(n4226), .Z(n4708) );
  CMXI2X1 U14249 ( .A0(n4706), .A1(n4708), .S(n3765), .Z(n4758) );
  CMXI2X1 U14250 ( .A0(n4934), .A1(n4611), .S(n3847), .Z(N122) );
  CMXI2X1 U14251 ( .A0(n4613), .A1(n4612), .S(n4215), .Z(n4672) );
  CMXI2X1 U14252 ( .A0(n4617), .A1(n4616), .S(n4219), .Z(n4674) );
  CMXI2X1 U14253 ( .A0(n4671), .A1(n4674), .S(n4226), .Z(n4712) );
  CMXI2X1 U14254 ( .A0(n4710), .A1(n4712), .S(n3762), .Z(n4760) );
  CMXI2X1 U14255 ( .A0(n4619), .A1(n4618), .S(n3247), .Z(n4673) );
  CMXI2X1 U14256 ( .A0(n4940), .A1(n4621), .S(n3848), .Z(N123) );
  CMXI2X1 U14257 ( .A0(n4623), .A1(n4622), .S(n4214), .Z(n4678) );
  CMXI2X1 U14258 ( .A0(n4627), .A1(n4626), .S(n4213), .Z(n4680) );
  CMXI2X1 U14259 ( .A0(n4714), .A1(n4716), .S(n3765), .Z(n4654) );
  CMXI2X1 U14260 ( .A0(n4629), .A1(n4628), .S(n4217), .Z(n4679) );
  CMXI2X1 U14261 ( .A0(n4679), .A1(n4681), .S(n4226), .Z(n4715) );
  CMXI2X1 U14262 ( .A0(n4946), .A1(n4631), .S(n3849), .Z(N124) );
  CMXI2X1 U14263 ( .A0(n4633), .A1(n4632), .S(n4214), .Z(n4684) );
  CMXI2X1 U14264 ( .A0(n4635), .A1(n4634), .S(n4219), .Z(n4683) );
  CMXI2X1 U14265 ( .A0(n4637), .A1(n4636), .S(n4218), .Z(n4686) );
  CMXI2X1 U14266 ( .A0(n4683), .A1(n4686), .S(n4227), .Z(n4720) );
  CMXI2X1 U14267 ( .A0(n4639), .A1(n4638), .S(n4215), .Z(n4685) );
  CMXI2X1 U14268 ( .A0(n4952), .A1(n4641), .S(n3850), .Z(N125) );
  CMXI2X1 U14269 ( .A0(n4644), .A1(n4643), .S(n4226), .Z(n4724) );
  CMXI2X1 U14270 ( .A0(n4722), .A1(n4724), .S(n3765), .Z(n4742) );
  CMXI2X1 U14271 ( .A0(n4646), .A1(n4645), .S(n4226), .Z(n4723) );
  CMXI2X1 U14272 ( .A0(n4958), .A1(n4647), .S(n3851), .Z(N126) );
  CMXI2X1 U14273 ( .A0(n4726), .A1(n4728), .S(n3766), .Z(n4764) );
  CMXI2X1 U14274 ( .A0(n4964), .A1(n4653), .S(n3852), .Z(N127) );
  CMX2X1 U14275 ( .A0(n4655), .A1(n4654), .S(n3205), .Z(n4884) );
  CMXI2X1 U14276 ( .A0(n4658), .A1(n4657), .S(n4226), .Z(n4732) );
  CMXI2X1 U14277 ( .A0(n4730), .A1(n4732), .S(n3763), .Z(n4768) );
  CMXI2X1 U14278 ( .A0(n4970), .A1(n4661), .S(n3853), .Z(N128) );
  CMXI2X1 U14279 ( .A0(n4664), .A1(n4663), .S(n4227), .Z(n4736) );
  CMXI2X1 U14280 ( .A0(n4734), .A1(n4736), .S(n3766), .Z(n4770) );
  CMXI2X1 U14281 ( .A0(n4666), .A1(n4665), .S(n4226), .Z(n4735) );
  CMXI2X1 U14282 ( .A0(n4976), .A1(n4667), .S(n3834), .Z(N129) );
  CMXI2X1 U14283 ( .A0(n4983), .A1(n4670), .S(n3843), .Z(N130) );
  CMXI2X1 U14284 ( .A0(n4672), .A1(n4671), .S(n4226), .Z(n4741) );
  CMXI2X1 U14285 ( .A0(n4674), .A1(n4673), .S(n4226), .Z(n4740) );
  CMXI2X1 U14286 ( .A0(n4740), .A1(n4739), .S(n3763), .Z(n4775) );
  CMXI2X1 U14287 ( .A0(n4990), .A1(n4676), .S(n3843), .Z(N131) );
  CMXI2X1 U14288 ( .A0(n4678), .A1(n4677), .S(n4226), .Z(n4746) );
  CMXI2X1 U14289 ( .A0(n4680), .A1(n4679), .S(n4226), .Z(n4745) );
  CMXI2X1 U14290 ( .A0(n4745), .A1(n4744), .S(n3766), .Z(n4777) );
  CMXI2X1 U14291 ( .A0(n4997), .A1(n4682), .S(n3844), .Z(N132) );
  CMXI2X1 U14292 ( .A0(n4684), .A1(n4683), .S(n4227), .Z(n4749) );
  CMXI2X1 U14293 ( .A0(n4686), .A1(n4685), .S(n4226), .Z(n4748) );
  CMXI2X1 U14294 ( .A0(n4748), .A1(n4747), .S(n3764), .Z(n4779) );
  CMXI2X1 U14295 ( .A0(n5004), .A1(n4688), .S(n3853), .Z(N133) );
  CMXI2X1 U14296 ( .A0(n4690), .A1(n4689), .S(n3764), .Z(n4781) );
  CMXI2X1 U14297 ( .A0(n5011), .A1(n4691), .S(n3845), .Z(N134) );
  CMXI2X1 U14298 ( .A0(n4694), .A1(n4693), .S(n3762), .Z(n4783) );
  CMXI2X1 U14299 ( .A0(n5018), .A1(n4695), .S(n3835), .Z(N135) );
  CMXI2X1 U14300 ( .A0(n4698), .A1(n4697), .S(n3764), .Z(n4786) );
  CMXI2X1 U14301 ( .A0(n5025), .A1(n4699), .S(n3836), .Z(N136) );
  CMXI2X1 U14302 ( .A0(n3699), .A1(n4701), .S(n3762), .Z(n4788) );
  CMXI2X1 U14303 ( .A0(n5032), .A1(n4703), .S(n3837), .Z(N137) );
  CMX2X1 U14304 ( .A0(n4705), .A1(n4704), .S(n3211), .Z(n4885) );
  CMXI2X1 U14305 ( .A0(n4708), .A1(n4707), .S(n3765), .Z(n4790) );
  CMXI2X1 U14306 ( .A0(n5039), .A1(n4709), .S(n3838), .Z(N138) );
  CMXI2X1 U14307 ( .A0(n4712), .A1(n4711), .S(n3765), .Z(n4792) );
  CMXI2X1 U14308 ( .A0(n5046), .A1(n4713), .S(n3835), .Z(N139) );
  CMXI2X1 U14309 ( .A0(n4716), .A1(n4715), .S(n3763), .Z(n4794) );
  CMXI2X1 U14310 ( .A0(n5054), .A1(n4717), .S(n3839), .Z(N140) );
  CMXI2X1 U14311 ( .A0(n3702), .A1(n4719), .S(n3703), .Z(n4796) );
  CMXI2X1 U14312 ( .A0(n5061), .A1(n4721), .S(n3840), .Z(N141) );
  CMXI2X1 U14313 ( .A0(n4724), .A1(n4723), .S(n3763), .Z(n4798) );
  CMXI2X1 U14314 ( .A0(n5068), .A1(n4725), .S(n3841), .Z(N142) );
  CMXI2X1 U14315 ( .A0(n4728), .A1(n4727), .S(n3766), .Z(n4800) );
  CMXI2X1 U14316 ( .A0(n5075), .A1(n4729), .S(n3842), .Z(N143) );
  CMXI2X1 U14317 ( .A0(n4732), .A1(n4731), .S(n3763), .Z(n4802) );
  CMXI2X1 U14318 ( .A0(n5082), .A1(n4733), .S(n3843), .Z(N144) );
  CMXI2X1 U14319 ( .A0(n4736), .A1(n4735), .S(n3766), .Z(n4804) );
  CMXI2X1 U14320 ( .A0(n5089), .A1(n4737), .S(n3844), .Z(N145) );
  CMXI2X1 U14321 ( .A0(n4741), .A1(n4740), .S(n3764), .Z(n4808) );
  CMX2X1 U14322 ( .A0(n4743), .A1(n4742), .S(n3209), .Z(n4886) );
  CMXI2X1 U14323 ( .A0(n4746), .A1(n4745), .S(n3762), .Z(n4810) );
  CMX2X1 U14324 ( .A0(n4809), .A1(n4810), .S(n3213), .Z(n4874) );
  CMXI2X1 U14325 ( .A0(n4749), .A1(n4748), .S(n3766), .Z(n4812) );
  CMX2X1 U14326 ( .A0(n4811), .A1(n4812), .S(n3201), .Z(n4875) );
  CMX2X1 U14327 ( .A0(n4751), .A1(n4750), .S(n3209), .Z(n4876) );
  CMX2X1 U14328 ( .A0(n4753), .A1(n4752), .S(n3199), .Z(n4877) );
  CMX2X1 U14329 ( .A0(n4759), .A1(n4758), .S(n3207), .Z(n4882) );
  CMX2X1 U14330 ( .A0(n4761), .A1(n4760), .S(n3211), .Z(n4883) );
  CMX2X1 U14331 ( .A0(n4765), .A1(n4764), .S(n3213), .Z(n4887) );
  CMX2X1 U14332 ( .A0(n4769), .A1(n4768), .S(n3209), .Z(n4888) );
  CMX2X1 U14333 ( .A0(n4771), .A1(n4770), .S(n3199), .Z(n4889) );
  CMX2X1 U14334 ( .A0(n4773), .A1(n4772), .S(n3211), .Z(n4890) );
  CMX2X1 U14335 ( .A0(n4775), .A1(n4774), .S(n3211), .Z(n4891) );
  CMX2X1 U14336 ( .A0(n4777), .A1(n4776), .S(n3203), .Z(n4893) );
  CMX2X1 U14337 ( .A0(n4779), .A1(n4778), .S(n3199), .Z(n4894) );
  CMX2X1 U14338 ( .A0(n4781), .A1(n4780), .S(n3209), .Z(n4895) );
  CMX2X1 U14339 ( .A0(n4783), .A1(n4782), .S(n3201), .Z(n4896) );
  CMX2X1 U14340 ( .A0(n4786), .A1(n4785), .S(n3213), .Z(n4897) );
  CMX2X1 U14341 ( .A0(n4788), .A1(n4787), .S(n3203), .Z(n4898) );
  CMX2X1 U14342 ( .A0(n4790), .A1(n4789), .S(n3211), .Z(n4899) );
  CMX2X1 U14343 ( .A0(n4792), .A1(n4791), .S(n3199), .Z(n4900) );
  CMX2X1 U14344 ( .A0(n4794), .A1(n4793), .S(n3215), .Z(n4901) );
  CMX2X1 U14345 ( .A0(n4796), .A1(n4795), .S(n3203), .Z(n4902) );
  CMX2X1 U14346 ( .A0(n3749), .A1(n4797), .S(n3215), .Z(n4904) );
  CMX2X1 U14347 ( .A0(n4800), .A1(n4799), .S(n3205), .Z(n4905) );
  CMX2X1 U14348 ( .A0(n4804), .A1(n4803), .S(n3199), .Z(n4907) );
  CMX2X1 U14349 ( .A0(n6486), .A1(n4909), .S(n3730), .Z(n5276) );
  CMX2X1 U14350 ( .A0(n6499), .A1(n4911), .S(n3726), .Z(n5287) );
  CMX2X1 U14351 ( .A0(n6512), .A1(n4914), .S(n3721), .Z(n5305) );
  CMXI2X1 U14352 ( .A0(n4814), .A1(n4813), .S(n3728), .Z(n5326) );
  CMXI2X1 U14353 ( .A0(n4816), .A1(n4815), .S(n3729), .Z(n5347) );
  CMXI2X1 U14354 ( .A0(n4818), .A1(n4817), .S(n3724), .Z(n5362) );
  CMXI2X1 U14355 ( .A0(n4820), .A1(n4819), .S(n3726), .Z(n5373) );
  CMXI2X1 U14356 ( .A0(n4822), .A1(n4821), .S(n3727), .Z(n5385) );
  CMXI2X1 U14357 ( .A0(n4824), .A1(n4823), .S(n3730), .Z(n5396) );
  CMXI2X1 U14358 ( .A0(n4827), .A1(n4826), .S(n3727), .Z(n5407) );
  CMXI2X1 U14359 ( .A0(n4829), .A1(n4828), .S(n3724), .Z(n5418) );
  CMXI2X1 U14360 ( .A0(n4831), .A1(n4830), .S(n3722), .Z(n5429) );
  CMXI2X1 U14361 ( .A0(n4833), .A1(n4832), .S(n3726), .Z(n5440) );
  CMXI2X1 U14362 ( .A0(n4835), .A1(n4834), .S(n3726), .Z(n5451) );
  CMXI2X1 U14363 ( .A0(n4837), .A1(n4836), .S(n3727), .Z(n5462) );
  CMXI2X1 U14364 ( .A0(n4839), .A1(n4838), .S(n3730), .Z(n5503) );
  CMXI2X1 U14365 ( .A0(n4841), .A1(n4840), .S(n3725), .Z(n5567) );
  CMXI2X1 U14366 ( .A0(n4843), .A1(n4842), .S(n3727), .Z(n5639) );
  CMXI2X1 U14367 ( .A0(n4845), .A1(n4844), .S(n3724), .Z(n5692) );
  CMXI2X1 U14368 ( .A0(n4848), .A1(n4847), .S(n3723), .Z(n5721) );
  CMXI2X1 U14369 ( .A0(n4850), .A1(n4849), .S(n3729), .Z(n5742) );
  CMXI2X1 U14370 ( .A0(n4852), .A1(n4851), .S(n3730), .Z(n5762) );
  CMXI2X1 U14371 ( .A0(n4854), .A1(n4853), .S(n3730), .Z(n5783) );
  CMXI2X1 U14372 ( .A0(n4856), .A1(n4855), .S(n3727), .Z(n5804) );
  CMXI2X1 U14373 ( .A0(n4858), .A1(n4857), .S(n3722), .Z(n5821) );
  CMXI2X1 U14374 ( .A0(n4860), .A1(n4859), .S(n3722), .Z(n5832) );
  CMXI2X1 U14375 ( .A0(n4862), .A1(n4861), .S(n3727), .Z(n5843) );
  CMXI2X1 U14376 ( .A0(n4864), .A1(n4863), .S(n3730), .Z(n5856) );
  CMXI2X1 U14377 ( .A0(n4866), .A1(n4865), .S(n3729), .Z(n5877) );
  CMXI2X1 U14378 ( .A0(n4869), .A1(n4868), .S(n3723), .Z(n5898) );
  CMXI2X1 U14379 ( .A0(n4871), .A1(n4870), .S(n3726), .Z(n5919) );
  CND2IX1 U14380 ( .B(n5189), .A(n3730), .Z(n5292) );
  CND2IX1 U14381 ( .B(n4909), .A(n3733), .Z(n6488) );
  CMXI2X1 U14382 ( .A0(n5292), .A1(n6488), .S(n3845), .Z(N243) );
  CMXI2X1 U14383 ( .A0(n4912), .A1(n4910), .S(n4211), .Z(n4916) );
  CND2IX1 U14384 ( .B(n5192), .A(n3724), .Z(n5294) );
  CND2IX1 U14385 ( .B(n4911), .A(n3733), .Z(n6501) );
  CMXI2X1 U14386 ( .A0(n5294), .A1(n6501), .S(n3846), .Z(N244) );
  CMXI2X1 U14387 ( .A0(n4915), .A1(n4912), .S(n4211), .Z(n4919) );
  CMXI2X1 U14388 ( .A0(n4919), .A1(n4913), .S(n3188), .Z(n4929) );
  CND2IX1 U14389 ( .B(n4914), .A(n3732), .Z(n6514) );
  CMXI2X1 U14390 ( .A0(n5296), .A1(n6514), .S(n3847), .Z(N245) );
  CMXI2X1 U14391 ( .A0(n4918), .A1(n4915), .S(n4209), .Z(n4924) );
  CMXI2X1 U14392 ( .A0(n4924), .A1(n4916), .S(n3188), .Z(n4933) );
  CND2IX1 U14393 ( .B(n5196), .A(n3727), .Z(n5298) );
  CMXI2X1 U14394 ( .A0(n5298), .A1(n4917), .S(n3848), .Z(N246) );
  CMXI2X1 U14395 ( .A0(n4923), .A1(n4918), .S(n4210), .Z(n4928) );
  CMXI2X1 U14396 ( .A0(n5300), .A1(n4921), .S(n3844), .Z(N247) );
  CMXI2X1 U14397 ( .A0(n4927), .A1(n4923), .S(n4203), .Z(n4932) );
  CMXI2X1 U14398 ( .A0(n4932), .A1(n4924), .S(n3194), .Z(n4944) );
  CMXI2X1 U14399 ( .A0(n4944), .A1(n4925), .S(n4217), .Z(n4969) );
  CMXI2X1 U14400 ( .A0(n5302), .A1(n4926), .S(n3846), .Z(N248) );
  CMXI2X1 U14401 ( .A0(n4931), .A1(n4927), .S(n4211), .Z(n4937) );
  CMXI2X1 U14402 ( .A0(n4937), .A1(n4928), .S(n3192), .Z(n4950) );
  CMXI2X1 U14403 ( .A0(n4950), .A1(n4929), .S(n3246), .Z(n4975) );
  CND2IX1 U14404 ( .B(n5202), .A(n3728), .Z(n5304) );
  CMXI2X1 U14405 ( .A0(n5304), .A1(n4930), .S(n3847), .Z(N249) );
  CMXI2X1 U14406 ( .A0(n4936), .A1(n4931), .S(n4208), .Z(n4943) );
  CMXI2X1 U14407 ( .A0(n4943), .A1(n4932), .S(n3188), .Z(n4956) );
  CMXI2X1 U14408 ( .A0(n4956), .A1(n4933), .S(n4215), .Z(n4982) );
  CND2IX1 U14409 ( .B(n5204), .A(n3722), .Z(n5307) );
  CMXI2X1 U14410 ( .A0(n5307), .A1(n4934), .S(n3834), .Z(N250) );
  CMXI2X1 U14411 ( .A0(n4942), .A1(n4936), .S(n4209), .Z(n4949) );
  CMXI2X1 U14412 ( .A0(n4949), .A1(n4937), .S(n3188), .Z(n4962) );
  CMXI2X1 U14413 ( .A0(n4962), .A1(n4938), .S(n4214), .Z(n4988) );
  CMXI2X1 U14414 ( .A0(n4988), .A1(n4939), .S(n4226), .Z(n5045) );
  CMXI2X1 U14415 ( .A0(n5309), .A1(n4940), .S(n3848), .Z(N251) );
  CMXI2X1 U14416 ( .A0(n4948), .A1(n4942), .S(n4206), .Z(n4955) );
  CMXI2X1 U14417 ( .A0(n4955), .A1(n4943), .S(n3188), .Z(n4968) );
  CMXI2X1 U14418 ( .A0(n4968), .A1(n4944), .S(n4216), .Z(n4995) );
  CMXI2X1 U14419 ( .A0(n4995), .A1(n4945), .S(n4223), .Z(n5053) );
  CMXI2X1 U14420 ( .A0(n5311), .A1(n4946), .S(n3849), .Z(N252) );
  CMXI2X1 U14421 ( .A0(n4954), .A1(n4948), .S(n4206), .Z(n4961) );
  CMXI2X1 U14422 ( .A0(n4961), .A1(n4949), .S(n3194), .Z(n4974) );
  CMXI2X1 U14423 ( .A0(n4974), .A1(n4950), .S(n4215), .Z(n5002) );
  CMXI2X1 U14424 ( .A0(n5002), .A1(n4951), .S(n4222), .Z(n5060) );
  CND2IX1 U14425 ( .B(n5210), .A(n3723), .Z(n5313) );
  CMXI2X1 U14426 ( .A0(n5313), .A1(n4952), .S(n3850), .Z(N253) );
  CMXI2X1 U14427 ( .A0(n4960), .A1(n4954), .S(n4208), .Z(n4967) );
  CMXI2X1 U14428 ( .A0(n4967), .A1(n4955), .S(n3192), .Z(n4981) );
  CMXI2X1 U14429 ( .A0(n4981), .A1(n4956), .S(n4213), .Z(n5009) );
  CMXI2X1 U14430 ( .A0(n5009), .A1(n4957), .S(n4225), .Z(n5067) );
  CND2IX1 U14431 ( .B(n5214), .A(n3723), .Z(n5315) );
  CMXI2X1 U14432 ( .A0(n5315), .A1(n4958), .S(n3851), .Z(N254) );
  CMXI2X1 U14433 ( .A0(n4966), .A1(n4960), .S(n4203), .Z(n4973) );
  CMXI2X1 U14434 ( .A0(n4973), .A1(n4961), .S(n3188), .Z(n4987) );
  CMXI2X1 U14435 ( .A0(n4987), .A1(n4962), .S(n4216), .Z(n5016) );
  CMXI2X1 U14436 ( .A0(n5016), .A1(n4963), .S(n4226), .Z(n5074) );
  CND2IX1 U14437 ( .B(n5216), .A(n3726), .Z(n5317) );
  CMXI2X1 U14438 ( .A0(n5317), .A1(n4964), .S(n3852), .Z(N255) );
  CMXI2X1 U14439 ( .A0(n4972), .A1(n4966), .S(n4211), .Z(n4980) );
  CMXI2X1 U14440 ( .A0(n4980), .A1(n4967), .S(n3194), .Z(n4994) );
  CMXI2X1 U14441 ( .A0(n5023), .A1(n4969), .S(n4226), .Z(n5081) );
  CND2IX1 U14442 ( .B(n5218), .A(n3729), .Z(n5319) );
  CMXI2X1 U14443 ( .A0(n5319), .A1(n4970), .S(n3836), .Z(N256) );
  CMXI2X1 U14444 ( .A0(n4979), .A1(n4972), .S(n4210), .Z(n4986) );
  CMXI2X1 U14445 ( .A0(n4986), .A1(n4973), .S(n3188), .Z(n5001) );
  CMXI2X1 U14446 ( .A0(n5001), .A1(n4974), .S(n4212), .Z(n5030) );
  CND2IX1 U14447 ( .B(n5220), .A(n3722), .Z(n5321) );
  CMXI2X1 U14448 ( .A0(n5321), .A1(n4976), .S(n3853), .Z(N257) );
  CMXI2X1 U14449 ( .A0(n4985), .A1(n4979), .S(n4206), .Z(n4993) );
  CMXI2X1 U14450 ( .A0(n4993), .A1(n4980), .S(n3192), .Z(n5008) );
  CMXI2X1 U14451 ( .A0(n5008), .A1(n4981), .S(n4218), .Z(n5037) );
  CMXI2X1 U14452 ( .A0(n5037), .A1(n4982), .S(n4226), .Z(n5095) );
  CND2IX1 U14453 ( .B(n5222), .A(n3729), .Z(n5323) );
  CMXI2X1 U14454 ( .A0(n5323), .A1(n4983), .S(n3834), .Z(N258) );
  CMXI2X1 U14455 ( .A0(n4992), .A1(n4985), .S(n4206), .Z(n5000) );
  CMXI2X1 U14456 ( .A0(n5000), .A1(n4986), .S(n3190), .Z(n5015) );
  CMXI2X1 U14457 ( .A0(n5015), .A1(n4987), .S(n4212), .Z(n5044) );
  CMXI2X1 U14458 ( .A0(n5044), .A1(n4988), .S(n4224), .Z(n5100) );
  CMXI2X1 U14459 ( .A0(n5100), .A1(n4989), .S(n3762), .Z(n5157) );
  CND2IX1 U14460 ( .B(n5224), .A(n3729), .Z(n5325) );
  CMXI2X1 U14461 ( .A0(n5325), .A1(n4990), .S(n3835), .Z(N259) );
  CMXI2X1 U14462 ( .A0(n4999), .A1(n4992), .S(n4205), .Z(n5007) );
  CMXI2X1 U14463 ( .A0(n5007), .A1(n4993), .S(n3188), .Z(n5022) );
  CMXI2X1 U14464 ( .A0(n5105), .A1(n4996), .S(n3240), .Z(n5159) );
  CND2IX1 U14465 ( .B(n5226), .A(n3724), .Z(n5328) );
  CMXI2X1 U14466 ( .A0(n5328), .A1(n4997), .S(n3836), .Z(N260) );
  CMXI2X1 U14467 ( .A0(n5006), .A1(n4999), .S(n4208), .Z(n5014) );
  CMXI2X1 U14468 ( .A0(n5014), .A1(n5000), .S(n3194), .Z(n5029) );
  CMXI2X1 U14469 ( .A0(n5029), .A1(n5001), .S(n4214), .Z(n5059) );
  CMXI2X1 U14470 ( .A0(n5059), .A1(n5002), .S(n4224), .Z(n5110) );
  CMXI2X1 U14471 ( .A0(n5110), .A1(n5003), .S(n3765), .Z(n5161) );
  CND2IX1 U14472 ( .B(n5228), .A(n3725), .Z(n5330) );
  CMXI2X1 U14473 ( .A0(n5330), .A1(n5004), .S(n3837), .Z(N261) );
  CMXI2X1 U14474 ( .A0(n5013), .A1(n5006), .S(n4209), .Z(n5021) );
  CMXI2X1 U14475 ( .A0(n5021), .A1(n5007), .S(n3188), .Z(n5036) );
  CMXI2X1 U14476 ( .A0(n5036), .A1(n5008), .S(n3247), .Z(n5066) );
  CMXI2X1 U14477 ( .A0(n5066), .A1(n5009), .S(n4226), .Z(n5115) );
  CMXI2X1 U14478 ( .A0(n5115), .A1(n5010), .S(n3765), .Z(n5163) );
  CND2IX1 U14479 ( .B(n5230), .A(n3725), .Z(n5332) );
  CMXI2X1 U14480 ( .A0(n5332), .A1(n5011), .S(n3838), .Z(N262) );
  CMXI2X1 U14481 ( .A0(n5020), .A1(n5013), .S(n4210), .Z(n5028) );
  CMXI2X1 U14482 ( .A0(n5028), .A1(n5014), .S(n3188), .Z(n5043) );
  CMXI2X1 U14483 ( .A0(n5043), .A1(n5015), .S(n4215), .Z(n5073) );
  CMXI2X1 U14484 ( .A0(n5073), .A1(n5016), .S(n4226), .Z(n5119) );
  CMXI2X1 U14485 ( .A0(n5119), .A1(n5017), .S(n3765), .Z(n5165) );
  CND2IX1 U14486 ( .B(n5232), .A(n3729), .Z(n5334) );
  CMXI2X1 U14487 ( .A0(n5334), .A1(n5018), .S(n3839), .Z(N263) );
  CMXI2X1 U14488 ( .A0(n5027), .A1(n5020), .S(n4203), .Z(n5035) );
  CMXI2X1 U14489 ( .A0(n5035), .A1(n5021), .S(n3188), .Z(n5051) );
  CMXI2X1 U14490 ( .A0(n5051), .A1(n5022), .S(n4218), .Z(n5080) );
  CMXI2X1 U14491 ( .A0(n5080), .A1(n5023), .S(n4224), .Z(n5123) );
  CMXI2X1 U14492 ( .A0(n5123), .A1(n5024), .S(n3763), .Z(n5167) );
  CND2IX1 U14493 ( .B(n5235), .A(n3723), .Z(n5336) );
  CMXI2X1 U14494 ( .A0(n5336), .A1(n5025), .S(n3840), .Z(N264) );
  CMXI2X1 U14495 ( .A0(n5034), .A1(n5027), .S(n4207), .Z(n5042) );
  CMXI2X1 U14496 ( .A0(n5042), .A1(n5028), .S(n3190), .Z(n5058) );
  CMXI2X1 U14497 ( .A0(n5058), .A1(n5029), .S(n3246), .Z(n5087) );
  CMXI2X1 U14498 ( .A0(n5127), .A1(n5031), .S(n3766), .Z(n5169) );
  CND2IX1 U14499 ( .B(n5237), .A(n3723), .Z(n5338) );
  CMXI2X1 U14500 ( .A0(n5338), .A1(n5032), .S(n3841), .Z(N265) );
  CMXI2X1 U14501 ( .A0(n5041), .A1(n5034), .S(n4205), .Z(n5050) );
  CMXI2X1 U14502 ( .A0(n5050), .A1(n5035), .S(n3192), .Z(n5065) );
  CMXI2X1 U14503 ( .A0(n5065), .A1(n5036), .S(n4215), .Z(n5094) );
  CMXI2X1 U14504 ( .A0(n3715), .A1(n5038), .S(n3764), .Z(n5172) );
  CND2IX1 U14505 ( .B(n5239), .A(n3728), .Z(n5340) );
  CMXI2X1 U14506 ( .A0(n5340), .A1(n5039), .S(n3842), .Z(N266) );
  CMXI2X1 U14507 ( .A0(n5049), .A1(n5041), .S(n4208), .Z(n5057) );
  CMXI2X1 U14508 ( .A0(n5057), .A1(n5042), .S(n3190), .Z(n5072) );
  CMXI2X1 U14509 ( .A0(n5072), .A1(n5043), .S(n4218), .Z(n5099) );
  CMXI2X1 U14510 ( .A0(n5099), .A1(n5044), .S(n4227), .Z(n5133) );
  CMXI2X1 U14511 ( .A0(n5133), .A1(n5045), .S(n3766), .Z(n5174) );
  CND2IX1 U14512 ( .B(n5241), .A(n3727), .Z(n5342) );
  CMXI2X1 U14513 ( .A0(n5342), .A1(n5046), .S(n3845), .Z(N267) );
  CMXI2X1 U14514 ( .A0(n5056), .A1(n5049), .S(n4211), .Z(n5064) );
  CMXI2X1 U14515 ( .A0(n5064), .A1(n5050), .S(n3190), .Z(n5079) );
  CMXI2X1 U14516 ( .A0(n5079), .A1(n5051), .S(n4215), .Z(n5104) );
  CMXI2X1 U14517 ( .A0(n5136), .A1(n5053), .S(n3762), .Z(n5176) );
  CND2IX1 U14518 ( .B(n5243), .A(n3722), .Z(n5344) );
  CMXI2X1 U14519 ( .A0(n5344), .A1(n5054), .S(n3849), .Z(N268) );
  CMXI2X1 U14520 ( .A0(n5063), .A1(n5056), .S(n4206), .Z(n5071) );
  CMXI2X1 U14521 ( .A0(n5071), .A1(n5057), .S(n3188), .Z(n5086) );
  CMXI2X1 U14522 ( .A0(n5086), .A1(n5058), .S(n4219), .Z(n5109) );
  CMXI2X1 U14523 ( .A0(n5109), .A1(n5059), .S(n4226), .Z(n5139) );
  CMXI2X1 U14524 ( .A0(n5139), .A1(n5060), .S(n3766), .Z(n5178) );
  CND2IX1 U14525 ( .B(n5245), .A(n3723), .Z(n5346) );
  CMXI2X1 U14526 ( .A0(n5346), .A1(n5061), .S(n3850), .Z(N269) );
  CMXI2X1 U14527 ( .A0(n5070), .A1(n5063), .S(n4204), .Z(n5078) );
  CMXI2X1 U14528 ( .A0(n5078), .A1(n5064), .S(n3190), .Z(n5093) );
  CMXI2X1 U14529 ( .A0(n5093), .A1(n5065), .S(n3246), .Z(n5114) );
  CMXI2X1 U14530 ( .A0(n5142), .A1(n5067), .S(n3764), .Z(n5180) );
  CND2IX1 U14531 ( .B(n5247), .A(n3726), .Z(n5349) );
  CMXI2X1 U14532 ( .A0(n5349), .A1(n5068), .S(n3835), .Z(N270) );
  CMXI2X1 U14533 ( .A0(n5077), .A1(n5070), .S(n4210), .Z(n5085) );
  CMXI2X1 U14534 ( .A0(n5085), .A1(n5071), .S(n3194), .Z(n5098) );
  CMXI2X1 U14535 ( .A0(n5098), .A1(n5072), .S(n4216), .Z(n5118) );
  CMXI2X1 U14536 ( .A0(n3719), .A1(n5074), .S(n3762), .Z(n5182) );
  CND2IX1 U14537 ( .B(n5249), .A(n3727), .Z(n5351) );
  CMXI2X1 U14538 ( .A0(n5351), .A1(n5075), .S(n3851), .Z(N271) );
  CMXI2X1 U14539 ( .A0(n5084), .A1(n5077), .S(n4207), .Z(n5092) );
  CMXI2X1 U14540 ( .A0(n5092), .A1(n5078), .S(n3194), .Z(n5103) );
  CMXI2X1 U14541 ( .A0(n5103), .A1(n5079), .S(n4215), .Z(n5122) );
  CMXI2X1 U14542 ( .A0(n5122), .A1(n5080), .S(n4226), .Z(n5149) );
  CMXI2X1 U14543 ( .A0(n5149), .A1(n5081), .S(n3766), .Z(n5184) );
  CND2IX1 U14544 ( .B(n5251), .A(n3726), .Z(n5353) );
  CMXI2X1 U14545 ( .A0(n5353), .A1(n5082), .S(n3843), .Z(N272) );
  CMXI2X1 U14546 ( .A0(n5091), .A1(n5084), .S(n4205), .Z(n5097) );
  CMXI2X1 U14547 ( .A0(n5097), .A1(n5085), .S(n3194), .Z(n5108) );
  CMXI2X1 U14548 ( .A0(n5108), .A1(n5086), .S(n4219), .Z(n5126) );
  CMXI2X1 U14549 ( .A0(n5126), .A1(n5087), .S(n4226), .Z(n5152) );
  CMXI2X1 U14550 ( .A0(n5152), .A1(n5088), .S(n3762), .Z(n5186) );
  CND2IX1 U14551 ( .B(n5253), .A(n3722), .Z(n5355) );
  CMXI2X1 U14552 ( .A0(n5355), .A1(n5089), .S(n3844), .Z(N273) );
  CMXI2X1 U14553 ( .A0(n5096), .A1(n5091), .S(n4206), .Z(n5102) );
  CMXI2X1 U14554 ( .A0(n5113), .A1(n5093), .S(n3246), .Z(n5129) );
  CMXI2X1 U14555 ( .A0(n5129), .A1(n5094), .S(n4226), .Z(n5154) );
  CMXI2X1 U14556 ( .A0(n5154), .A1(n5095), .S(n3763), .Z(n5187) );
  CMXI2X1 U14557 ( .A0(n5107), .A1(n5097), .S(n3190), .Z(n5117) );
  CMXI2X1 U14558 ( .A0(n5117), .A1(n5098), .S(n4219), .Z(n5132) );
  CMXI2X1 U14559 ( .A0(n5132), .A1(n5099), .S(n4226), .Z(n5156) );
  CMXI2X1 U14560 ( .A0(n5156), .A1(n5100), .S(n3763), .Z(n5188) );
  CMXI2X1 U14561 ( .A0(n5121), .A1(n5103), .S(n4213), .Z(n5135) );
  CMXI2X1 U14562 ( .A0(n5135), .A1(n5104), .S(n4222), .Z(n5158) );
  CMXI2X1 U14563 ( .A0(n5158), .A1(n3742), .S(n3765), .Z(n5191) );
  CMXI2X1 U14564 ( .A0(n5125), .A1(n5108), .S(n4217), .Z(n5138) );
  CMXI2X1 U14565 ( .A0(n5138), .A1(n5109), .S(n4223), .Z(n5160) );
  CMXI2X1 U14566 ( .A0(n5160), .A1(n5110), .S(n3766), .Z(n5193) );
  CMXI2X1 U14567 ( .A0(n5141), .A1(n5114), .S(n4226), .Z(n5162) );
  CMXI2X1 U14568 ( .A0(n5162), .A1(n5115), .S(n3766), .Z(n5195) );
  CMXI2X1 U14569 ( .A0(n5144), .A1(n5118), .S(n4226), .Z(n5164) );
  CMXI2X1 U14570 ( .A0(n5164), .A1(n5119), .S(n3762), .Z(n5197) );
  CMX2X1 U14571 ( .A0(n5120), .A1(n5197), .S(n3207), .Z(n5260) );
  CMXI2X1 U14572 ( .A0(n5148), .A1(n5122), .S(n4223), .Z(n5166) );
  CMXI2X1 U14573 ( .A0(n5166), .A1(n5123), .S(n3763), .Z(n5199) );
  CMXI2X1 U14574 ( .A0(n5151), .A1(n5126), .S(n4222), .Z(n5168) );
  CMXI2X1 U14575 ( .A0(n5168), .A1(n5127), .S(n3764), .Z(n5201) );
  CMX2X1 U14576 ( .A0(n5128), .A1(n5201), .S(n3211), .Z(n5262) );
  CMXI2X1 U14577 ( .A0(n5171), .A1(n5130), .S(n3766), .Z(n5203) );
  CMXI2X1 U14578 ( .A0(n5173), .A1(n5133), .S(n3763), .Z(n5205) );
  CMXI2X1 U14579 ( .A0(n5175), .A1(n5136), .S(n3762), .Z(n5207) );
  CMXI2X1 U14580 ( .A0(n5177), .A1(n5139), .S(n3765), .Z(n5209) );
  CMX2X1 U14581 ( .A0(n5140), .A1(n5209), .S(n3201), .Z(n5267) );
  CMXI2X1 U14582 ( .A0(n5179), .A1(n5142), .S(n3764), .Z(n5213) );
  CMXI2X1 U14583 ( .A0(n3717), .A1(n5145), .S(n3718), .Z(n5215) );
  CMXI2X1 U14584 ( .A0(n5183), .A1(n5149), .S(n3766), .Z(n5217) );
  CMXI2X1 U14585 ( .A0(n5185), .A1(n5152), .S(n3765), .Z(n5219) );
  CMX2X1 U14586 ( .A0(n5153), .A1(n5219), .S(n3213), .Z(n5271) );
  CMX2X1 U14587 ( .A0(n5155), .A1(n5221), .S(n3211), .Z(n5272) );
  CMX2X1 U14588 ( .A0(n5157), .A1(n5223), .S(n3205), .Z(n5273) );
  CMX2X1 U14589 ( .A0(n5159), .A1(n5225), .S(n3215), .Z(n5274) );
  CMX2X1 U14590 ( .A0(n5161), .A1(n5227), .S(n3213), .Z(n5275) );
  CMX2X1 U14591 ( .A0(n5163), .A1(n5229), .S(n3203), .Z(n5277) );
  CMX2X1 U14592 ( .A0(n5165), .A1(n5231), .S(n3203), .Z(n5278) );
  CMX2X1 U14593 ( .A0(n5167), .A1(n5234), .S(n3199), .Z(n5279) );
  CMX2X1 U14594 ( .A0(n5169), .A1(n5236), .S(n3215), .Z(n5280) );
  CMX2X1 U14595 ( .A0(n5172), .A1(n5238), .S(n3207), .Z(n5281) );
  CMX2X1 U14596 ( .A0(n5174), .A1(n5240), .S(n3211), .Z(n5282) );
  CMX2X1 U14597 ( .A0(n5176), .A1(n5242), .S(n3199), .Z(n5283) );
  CMX2X1 U14598 ( .A0(n5178), .A1(n5244), .S(n3205), .Z(n5284) );
  CMX2X1 U14599 ( .A0(n5180), .A1(n5246), .S(n3203), .Z(n5285) );
  CMX2X1 U14600 ( .A0(n5184), .A1(n5250), .S(n3211), .Z(n5288) );
  CMX2X1 U14601 ( .A0(n5186), .A1(n5252), .S(n3201), .Z(n5289) );
  CMX2X1 U14602 ( .A0(n5189), .A1(n5291), .S(n3726), .Z(n5393) );
  CMX2X1 U14603 ( .A0(n5192), .A1(n5293), .S(n3727), .Z(n5394) );
  CMX2X1 U14604 ( .A0(n5194), .A1(n5295), .S(n3721), .Z(n5395) );
  CMX2X1 U14605 ( .A0(n5196), .A1(n5297), .S(n3728), .Z(n5397) );
  CMX2X1 U14606 ( .A0(n5198), .A1(n5299), .S(n3729), .Z(n5398) );
  CMX2X1 U14607 ( .A0(n5200), .A1(n5301), .S(n3721), .Z(n5399) );
  CMX2X1 U14608 ( .A0(n5202), .A1(n5303), .S(n3725), .Z(n5400) );
  CMX2X1 U14609 ( .A0(n5204), .A1(n5306), .S(n3722), .Z(n5401) );
  CMX2X1 U14610 ( .A0(n5206), .A1(n5308), .S(n3729), .Z(n5402) );
  CMX2X1 U14611 ( .A0(n5208), .A1(n5310), .S(n3722), .Z(n5403) );
  CMX2X1 U14612 ( .A0(n5210), .A1(n5312), .S(n3729), .Z(n5404) );
  CMX2X1 U14613 ( .A0(n5214), .A1(n5314), .S(n3725), .Z(n5405) );
  CMX2X1 U14614 ( .A0(n5216), .A1(n5316), .S(n3730), .Z(n5406) );
  CMX2X1 U14615 ( .A0(n5218), .A1(n5318), .S(n3721), .Z(n5408) );
  CMX2X1 U14616 ( .A0(n5220), .A1(n5320), .S(n3725), .Z(n5409) );
  CMX2X1 U14617 ( .A0(n5222), .A1(n5322), .S(n3724), .Z(n5410) );
  CMX2X1 U14618 ( .A0(n5224), .A1(n5324), .S(n3730), .Z(n5411) );
  CMX2X1 U14619 ( .A0(n5226), .A1(n5327), .S(n3730), .Z(n5412) );
  CMX2X1 U14620 ( .A0(n5228), .A1(n5329), .S(n3728), .Z(n5413) );
  CMX2X1 U14621 ( .A0(n5230), .A1(n5331), .S(n3727), .Z(n5414) );
  CMX2X1 U14622 ( .A0(n5232), .A1(n5333), .S(n3723), .Z(n5415) );
  CMX2X1 U14623 ( .A0(n5235), .A1(n5335), .S(n3726), .Z(n5416) );
  CMX2X1 U14624 ( .A0(n5237), .A1(n5337), .S(n3727), .Z(n5417) );
  CMX2X1 U14625 ( .A0(n5239), .A1(n5339), .S(n3722), .Z(n5419) );
  CMX2X1 U14626 ( .A0(n5241), .A1(n5341), .S(n3729), .Z(n5420) );
  CMX2X1 U14627 ( .A0(n5243), .A1(n5343), .S(n3722), .Z(n5421) );
  CMX2X1 U14628 ( .A0(n5245), .A1(n5345), .S(n3726), .Z(n5422) );
  CMX2X1 U14629 ( .A0(n5247), .A1(n5348), .S(n3725), .Z(n5423) );
  CMX2X1 U14630 ( .A0(n5251), .A1(n5352), .S(n3724), .Z(n5425) );
  CND2IX1 U14631 ( .B(n5291), .A(n3732), .Z(n5465) );
  CMXI2X1 U14632 ( .A0(n5465), .A1(n5292), .S(n3845), .Z(N371) );
  CND2IX1 U14633 ( .B(n5293), .A(n3739), .Z(n5468) );
  CMXI2X1 U14634 ( .A0(n5468), .A1(n5294), .S(n3846), .Z(N372) );
  CND2IX1 U14635 ( .B(n5295), .A(n3736), .Z(n5472) );
  CMXI2X1 U14636 ( .A0(n5472), .A1(n5296), .S(n3837), .Z(N373) );
  CND2IX1 U14637 ( .B(n5297), .A(n3735), .Z(n5476) );
  CMXI2X1 U14638 ( .A0(n5476), .A1(n5298), .S(n3847), .Z(N374) );
  CND2IX1 U14639 ( .B(n5299), .A(n3735), .Z(n5481) );
  CMXI2X1 U14640 ( .A0(n5481), .A1(n5300), .S(n3848), .Z(N375) );
  CND2IX1 U14641 ( .B(n5301), .A(n3734), .Z(n5486) );
  CMXI2X1 U14642 ( .A0(n5486), .A1(n5302), .S(n3849), .Z(N376) );
  CND2IX1 U14643 ( .B(n5303), .A(n3740), .Z(n5491) );
  CMXI2X1 U14644 ( .A0(n5491), .A1(n5304), .S(n3850), .Z(N377) );
  CND2IX1 U14645 ( .B(n5306), .A(n3732), .Z(n5496) );
  CMXI2X1 U14646 ( .A0(n5496), .A1(n5307), .S(n3851), .Z(N378) );
  CND2IX1 U14647 ( .B(n5308), .A(n3732), .Z(n5502) );
  CMXI2X1 U14648 ( .A0(n5502), .A1(n5309), .S(n3852), .Z(N379) );
  CND2IX1 U14649 ( .B(n5310), .A(n3734), .Z(n5509) );
  CMXI2X1 U14650 ( .A0(n5509), .A1(n5311), .S(n3853), .Z(N380) );
  CND2IX1 U14651 ( .B(n5312), .A(n3738), .Z(n5515) );
  CMXI2X1 U14652 ( .A0(n5515), .A1(n5313), .S(n3834), .Z(N381) );
  CND2IX1 U14653 ( .B(n5314), .A(n3740), .Z(n5521) );
  CMXI2X1 U14654 ( .A0(n5521), .A1(n5315), .S(n3835), .Z(N382) );
  CND2IX1 U14655 ( .B(n5316), .A(n3738), .Z(n5527) );
  CMXI2X1 U14656 ( .A0(n5527), .A1(n5317), .S(n3836), .Z(N383) );
  CND2IX1 U14657 ( .B(n5318), .A(n3736), .Z(n5533) );
  CMXI2X1 U14658 ( .A0(n5533), .A1(n5319), .S(n3846), .Z(N384) );
  CND2IX1 U14659 ( .B(n5320), .A(n3733), .Z(n5539) );
  CMXI2X1 U14660 ( .A0(n5539), .A1(n5321), .S(n3852), .Z(N385) );
  CND2IX1 U14661 ( .B(n5322), .A(n3734), .Z(n5545) );
  CMXI2X1 U14662 ( .A0(n5545), .A1(n5323), .S(n3853), .Z(N386) );
  CND2IX1 U14663 ( .B(n5324), .A(n3735), .Z(n5552) );
  CMXI2X1 U14664 ( .A0(n5552), .A1(n5325), .S(n3836), .Z(N387) );
  CND2IX1 U14665 ( .B(n5327), .A(n3736), .Z(n5559) );
  CMXI2X1 U14666 ( .A0(n5559), .A1(n5328), .S(n3834), .Z(N388) );
  CND2IX1 U14667 ( .B(n5329), .A(n3737), .Z(n5566) );
  CMXI2X1 U14668 ( .A0(n5566), .A1(n5330), .S(n3837), .Z(N389) );
  CND2IX1 U14669 ( .B(n5331), .A(n3738), .Z(n5575) );
  CMXI2X1 U14670 ( .A0(n5575), .A1(n5332), .S(n3838), .Z(N390) );
  CND2IX1 U14671 ( .B(n5333), .A(n3736), .Z(n5582) );
  CMXI2X1 U14672 ( .A0(n5582), .A1(n5334), .S(n3839), .Z(N391) );
  CND2IX1 U14673 ( .B(n5335), .A(n3737), .Z(n5589) );
  CMXI2X1 U14674 ( .A0(n5589), .A1(n5336), .S(n3840), .Z(N392) );
  CND2IX1 U14675 ( .B(n5337), .A(n3738), .Z(n5596) );
  CMXI2X1 U14676 ( .A0(n5596), .A1(n5338), .S(n3838), .Z(N393) );
  CND2IX1 U14677 ( .B(n5339), .A(n3739), .Z(n5603) );
  CMXI2X1 U14678 ( .A0(n5603), .A1(n5340), .S(n3841), .Z(N394) );
  CMXI2X1 U14679 ( .A0(n5610), .A1(n5342), .S(n3842), .Z(N395) );
  CMXI2X1 U14680 ( .A0(n5617), .A1(n5344), .S(n3843), .Z(N396) );
  CMXI2X1 U14681 ( .A0(n5624), .A1(n5346), .S(n3844), .Z(N397) );
  CMXI2X1 U14682 ( .A0(n5631), .A1(n5349), .S(n3845), .Z(N398) );
  CMXI2X1 U14683 ( .A0(n5638), .A1(n5351), .S(n3846), .Z(N399) );
  CMXI2X1 U14684 ( .A0(n5646), .A1(n5353), .S(n3847), .Z(N400) );
  CMXI2X1 U14685 ( .A0(n5653), .A1(n5355), .S(n3848), .Z(N401) );
  CND2IX1 U14686 ( .B(n5753), .A(n3729), .Z(n5855) );
  CMXI2X1 U14687 ( .A0(n5855), .A1(n5465), .S(n3849), .Z(N499) );
  CMXI2X1 U14688 ( .A0(n5470), .A1(n5467), .S(n4206), .Z(n5475) );
  CND2IX1 U14689 ( .B(n5755), .A(n3728), .Z(n5858) );
  CMXI2X1 U14690 ( .A0(n5858), .A1(n5468), .S(n3850), .Z(N500) );
  CMXI2X1 U14691 ( .A0(n5474), .A1(n5470), .S(n4207), .Z(n5479) );
  CMXI2X1 U14692 ( .A0(n5479), .A1(n5471), .S(n3188), .Z(n5490) );
  CMXI2X1 U14693 ( .A0(n5860), .A1(n5472), .S(n3847), .Z(N501) );
  CMXI2X1 U14694 ( .A0(n5478), .A1(n5474), .S(n4209), .Z(n5484) );
  CMXI2X1 U14695 ( .A0(n5484), .A1(n5475), .S(n3192), .Z(n5495) );
  CND2IX1 U14696 ( .B(n5759), .A(n3730), .Z(n5862) );
  CMXI2X1 U14697 ( .A0(n5862), .A1(n5476), .S(n3835), .Z(N502) );
  CMXI2X1 U14698 ( .A0(n5483), .A1(n5478), .S(n4209), .Z(n5489) );
  CMXI2X1 U14699 ( .A0(n5489), .A1(n5479), .S(n3190), .Z(n5500) );
  CMXI2X1 U14700 ( .A0(n5500), .A1(n5480), .S(n4217), .Z(n5526) );
  CMXI2X1 U14701 ( .A0(n5864), .A1(n5481), .S(n3836), .Z(N503) );
  CMXI2X1 U14702 ( .A0(n5488), .A1(n5483), .S(n4204), .Z(n5494) );
  CMXI2X1 U14703 ( .A0(n5494), .A1(n5484), .S(n3190), .Z(n5507) );
  CMXI2X1 U14704 ( .A0(n5507), .A1(n5485), .S(n4213), .Z(n5532) );
  CMXI2X1 U14705 ( .A0(n5866), .A1(n5486), .S(n3837), .Z(N504) );
  CMXI2X1 U14706 ( .A0(n5493), .A1(n5488), .S(n4211), .Z(n5499) );
  CMXI2X1 U14707 ( .A0(n5499), .A1(n5489), .S(n3192), .Z(n5513) );
  CMXI2X1 U14708 ( .A0(n5513), .A1(n5490), .S(n4217), .Z(n5538) );
  CMXI2X1 U14709 ( .A0(n5868), .A1(n5491), .S(n3837), .Z(N505) );
  CMXI2X1 U14710 ( .A0(n5498), .A1(n5493), .S(n4205), .Z(n5506) );
  CMXI2X1 U14711 ( .A0(n5506), .A1(n5494), .S(n3192), .Z(n5519) );
  CMXI2X1 U14712 ( .A0(n5519), .A1(n5495), .S(n4212), .Z(n5544) );
  CND2IX1 U14713 ( .B(n5768), .A(n3726), .Z(n5870) );
  CMXI2X1 U14714 ( .A0(n5870), .A1(n5496), .S(n3851), .Z(N506) );
  CMXI2X1 U14715 ( .A0(n5505), .A1(n5498), .S(n4209), .Z(n5512) );
  CMXI2X1 U14716 ( .A0(n5512), .A1(n5499), .S(n3190), .Z(n5525) );
  CMXI2X1 U14717 ( .A0(n5525), .A1(n5500), .S(n4218), .Z(n5550) );
  CMXI2X1 U14718 ( .A0(n5550), .A1(n5501), .S(n4225), .Z(n5609) );
  CMXI2X1 U14719 ( .A0(n5872), .A1(n5502), .S(n3852), .Z(N507) );
  CMXI2X1 U14720 ( .A0(n5511), .A1(n5505), .S(n4211), .Z(n5518) );
  CMXI2X1 U14721 ( .A0(n5518), .A1(n5506), .S(n3194), .Z(n5531) );
  CMXI2X1 U14722 ( .A0(n5531), .A1(n5507), .S(n4217), .Z(n5557) );
  CMXI2X1 U14723 ( .A0(n5557), .A1(n5508), .S(n4226), .Z(n5616) );
  CMXI2X1 U14724 ( .A0(n5874), .A1(n5509), .S(n3853), .Z(N508) );
  CMXI2X1 U14725 ( .A0(n5517), .A1(n5511), .S(n4209), .Z(n5524) );
  CMXI2X1 U14726 ( .A0(n5524), .A1(n5512), .S(n3188), .Z(n5537) );
  CMXI2X1 U14727 ( .A0(n5537), .A1(n5513), .S(n3247), .Z(n5564) );
  CMXI2X1 U14728 ( .A0(n5564), .A1(n5514), .S(n4221), .Z(n5623) );
  CMXI2X1 U14729 ( .A0(n5876), .A1(n5515), .S(n3834), .Z(N509) );
  CMXI2X1 U14730 ( .A0(n5523), .A1(n5517), .S(n4207), .Z(n5530) );
  CMXI2X1 U14731 ( .A0(n5530), .A1(n5518), .S(n3194), .Z(n5543) );
  CMXI2X1 U14732 ( .A0(n5543), .A1(n5519), .S(n4212), .Z(n5573) );
  CMXI2X1 U14733 ( .A0(n5573), .A1(n5520), .S(n4224), .Z(n5630) );
  CMXI2X1 U14734 ( .A0(n5879), .A1(n5521), .S(n3839), .Z(N510) );
  CMXI2X1 U14735 ( .A0(n5529), .A1(n5523), .S(n4203), .Z(n5536) );
  CMXI2X1 U14736 ( .A0(n5536), .A1(n5524), .S(n3190), .Z(n5549) );
  CMXI2X1 U14737 ( .A0(n5549), .A1(n5525), .S(n4214), .Z(n5580) );
  CMXI2X1 U14738 ( .A0(n5580), .A1(n5526), .S(n4222), .Z(n5637) );
  CMXI2X1 U14739 ( .A0(n5881), .A1(n5527), .S(n3835), .Z(N511) );
  CMXI2X1 U14740 ( .A0(n5535), .A1(n5529), .S(n4210), .Z(n5542) );
  CMXI2X1 U14741 ( .A0(n5542), .A1(n5530), .S(n3192), .Z(n5556) );
  CMXI2X1 U14742 ( .A0(n5556), .A1(n5531), .S(n4215), .Z(n5587) );
  CMXI2X1 U14743 ( .A0(n5587), .A1(n5532), .S(n4226), .Z(n5645) );
  CMXI2X1 U14744 ( .A0(n5883), .A1(n5533), .S(n3836), .Z(N512) );
  CMXI2X1 U14745 ( .A0(n5541), .A1(n5535), .S(n4205), .Z(n5548) );
  CMXI2X1 U14746 ( .A0(n5548), .A1(n5536), .S(n3190), .Z(n5563) );
  CMXI2X1 U14747 ( .A0(n5563), .A1(n5537), .S(n4216), .Z(n5594) );
  CMXI2X1 U14748 ( .A0(n5594), .A1(n5538), .S(n4226), .Z(n5652) );
  CND2IX1 U14749 ( .B(n5782), .A(n3723), .Z(n5885) );
  CMXI2X1 U14750 ( .A0(n5885), .A1(n5539), .S(n3837), .Z(N513) );
  CMXI2X1 U14751 ( .A0(n5547), .A1(n5541), .S(n4208), .Z(n5555) );
  CMXI2X1 U14752 ( .A0(n5555), .A1(n5542), .S(n3192), .Z(n5572) );
  CMXI2X1 U14753 ( .A0(n5572), .A1(n5543), .S(n4220), .Z(n5601) );
  CMXI2X1 U14754 ( .A0(n5601), .A1(n5544), .S(n4226), .Z(n5659) );
  CND2IX1 U14755 ( .B(n5785), .A(n3727), .Z(n5887) );
  CMXI2X1 U14756 ( .A0(n5887), .A1(n5545), .S(n3838), .Z(N514) );
  CMXI2X1 U14757 ( .A0(n5554), .A1(n5547), .S(n4204), .Z(n5562) );
  CMXI2X1 U14758 ( .A0(n5562), .A1(n5548), .S(n3194), .Z(n5579) );
  CMXI2X1 U14759 ( .A0(n5579), .A1(n5549), .S(n4218), .Z(n5608) );
  CMXI2X1 U14760 ( .A0(n5608), .A1(n5550), .S(n4227), .Z(n5664) );
  CMXI2X1 U14761 ( .A0(n5664), .A1(n5551), .S(n3764), .Z(n5720) );
  CND2IX1 U14762 ( .B(n5787), .A(n3722), .Z(n5889) );
  CMXI2X1 U14763 ( .A0(n5889), .A1(n5552), .S(n3839), .Z(N515) );
  CMXI2X1 U14764 ( .A0(n5561), .A1(n5554), .S(n4203), .Z(n5571) );
  CMXI2X1 U14765 ( .A0(n5571), .A1(n5555), .S(n3194), .Z(n5586) );
  CMXI2X1 U14766 ( .A0(n5586), .A1(n5556), .S(n3246), .Z(n5615) );
  CMXI2X1 U14767 ( .A0(n5615), .A1(n5557), .S(n4227), .Z(n5669) );
  CMXI2X1 U14768 ( .A0(n5669), .A1(n5558), .S(n3762), .Z(n5723) );
  CMXI2X1 U14769 ( .A0(n5891), .A1(n5559), .S(n3840), .Z(N516) );
  CMXI2X1 U14770 ( .A0(n5570), .A1(n5561), .S(n4204), .Z(n5578) );
  CMXI2X1 U14771 ( .A0(n5578), .A1(n5562), .S(n3188), .Z(n5593) );
  CMXI2X1 U14772 ( .A0(n5593), .A1(n5563), .S(n4217), .Z(n5622) );
  CMXI2X1 U14773 ( .A0(n5622), .A1(n5564), .S(n4227), .Z(n5674) );
  CMXI2X1 U14774 ( .A0(n5674), .A1(n5565), .S(n3764), .Z(n5725) );
  CND2IX1 U14775 ( .B(n5791), .A(n3724), .Z(n5893) );
  CMXI2X1 U14776 ( .A0(n5893), .A1(n5566), .S(n3841), .Z(N517) );
  CMXI2X1 U14777 ( .A0(n5577), .A1(n5570), .S(n4208), .Z(n5585) );
  CMXI2X1 U14778 ( .A0(n5585), .A1(n5571), .S(n3192), .Z(n5600) );
  CMXI2X1 U14779 ( .A0(n5600), .A1(n5572), .S(n4215), .Z(n5629) );
  CMXI2X1 U14780 ( .A0(n5629), .A1(n5573), .S(n4227), .Z(n5678) );
  CMXI2X1 U14781 ( .A0(n5678), .A1(n5574), .S(n3766), .Z(n5727) );
  CND2IX1 U14782 ( .B(n5793), .A(n3730), .Z(n5895) );
  CMXI2X1 U14783 ( .A0(n5895), .A1(n5575), .S(n3842), .Z(N518) );
  CMXI2X1 U14784 ( .A0(n5584), .A1(n5577), .S(n4210), .Z(n5592) );
  CMXI2X1 U14785 ( .A0(n5592), .A1(n5578), .S(n3188), .Z(n5607) );
  CMXI2X1 U14786 ( .A0(n5607), .A1(n5579), .S(n4219), .Z(n5636) );
  CMXI2X1 U14787 ( .A0(n5636), .A1(n5580), .S(n4227), .Z(n5682) );
  CMXI2X1 U14788 ( .A0(n5682), .A1(n5581), .S(n3764), .Z(n5729) );
  CND2IX1 U14789 ( .B(n5795), .A(n3725), .Z(n5897) );
  CMXI2X1 U14790 ( .A0(n5897), .A1(n5582), .S(n3843), .Z(N519) );
  CMXI2X1 U14791 ( .A0(n5591), .A1(n5584), .S(n4203), .Z(n5599) );
  CMXI2X1 U14792 ( .A0(n5599), .A1(n5585), .S(n3194), .Z(n5614) );
  CMXI2X1 U14793 ( .A0(n5614), .A1(n5586), .S(n4216), .Z(n5644) );
  CMXI2X1 U14794 ( .A0(n5644), .A1(n5587), .S(n4227), .Z(n5686) );
  CMXI2X1 U14795 ( .A0(n5686), .A1(n5588), .S(n3763), .Z(n5731) );
  CND2IX1 U14796 ( .B(n5797), .A(n3728), .Z(n5900) );
  CMXI2X1 U14797 ( .A0(n5900), .A1(n5589), .S(n3844), .Z(N520) );
  CMXI2X1 U14798 ( .A0(n5598), .A1(n5591), .S(n4211), .Z(n5606) );
  CMXI2X1 U14799 ( .A0(n5606), .A1(n5592), .S(n3190), .Z(n5621) );
  CMXI2X1 U14800 ( .A0(n5621), .A1(n5593), .S(n4219), .Z(n5651) );
  CMXI2X1 U14801 ( .A0(n5651), .A1(n5594), .S(n4227), .Z(n5690) );
  CMXI2X1 U14802 ( .A0(n5690), .A1(n5595), .S(n3766), .Z(n5733) );
  CND2IX1 U14803 ( .B(n5799), .A(n3727), .Z(n5902) );
  CMXI2X1 U14804 ( .A0(n5902), .A1(n5596), .S(n3848), .Z(N521) );
  CMXI2X1 U14805 ( .A0(n5605), .A1(n5598), .S(n4204), .Z(n5613) );
  CMXI2X1 U14806 ( .A0(n5613), .A1(n5599), .S(n3192), .Z(n5628) );
  CMXI2X1 U14807 ( .A0(n5628), .A1(n5600), .S(n4213), .Z(n5658) );
  CMXI2X1 U14808 ( .A0(n5658), .A1(n5601), .S(n4227), .Z(n5694) );
  CMXI2X1 U14809 ( .A0(n5694), .A1(n5602), .S(n3763), .Z(n5735) );
  CND2IX1 U14810 ( .B(n5801), .A(n3722), .Z(n5904) );
  CMXI2X1 U14811 ( .A0(n5904), .A1(n5603), .S(n3838), .Z(N522) );
  CMXI2X1 U14812 ( .A0(n5612), .A1(n5605), .S(n4205), .Z(n5620) );
  CMXI2X1 U14813 ( .A0(n5620), .A1(n5606), .S(n3194), .Z(n5635) );
  CMXI2X1 U14814 ( .A0(n5635), .A1(n5607), .S(n4218), .Z(n5663) );
  CMXI2X1 U14815 ( .A0(n5663), .A1(n5608), .S(n4227), .Z(n5697) );
  CMXI2X1 U14816 ( .A0(n5697), .A1(n5609), .S(n3763), .Z(n5737) );
  CND2IX1 U14817 ( .B(n5803), .A(n3724), .Z(n5906) );
  CMXI2X1 U14818 ( .A0(n5906), .A1(n5610), .S(n3839), .Z(N523) );
  CMXI2X1 U14819 ( .A0(n5619), .A1(n5612), .S(n4210), .Z(n5627) );
  CMXI2X1 U14820 ( .A0(n5627), .A1(n5613), .S(n3192), .Z(n5643) );
  CMXI2X1 U14821 ( .A0(n5643), .A1(n5614), .S(n4218), .Z(n5668) );
  CMXI2X1 U14822 ( .A0(n5668), .A1(n5615), .S(n4227), .Z(n5700) );
  CMXI2X1 U14823 ( .A0(n5700), .A1(n5616), .S(n3766), .Z(n5739) );
  CND2IX1 U14824 ( .B(n5806), .A(n3722), .Z(n5908) );
  CMXI2X1 U14825 ( .A0(n5908), .A1(n5617), .S(n3838), .Z(N524) );
  CMXI2X1 U14826 ( .A0(n5626), .A1(n5619), .S(n4206), .Z(n5634) );
  CMXI2X1 U14827 ( .A0(n5634), .A1(n5620), .S(n3192), .Z(n5650) );
  CMXI2X1 U14828 ( .A0(n5650), .A1(n5621), .S(n4217), .Z(n5673) );
  CMXI2X1 U14829 ( .A0(n5673), .A1(n5622), .S(n4224), .Z(n5703) );
  CMXI2X1 U14830 ( .A0(n5703), .A1(n5623), .S(n3765), .Z(n5741) );
  CND2IX1 U14831 ( .B(n5808), .A(n3725), .Z(n5910) );
  CMXI2X1 U14832 ( .A0(n5910), .A1(n5624), .S(n3840), .Z(N525) );
  CMXI2X1 U14833 ( .A0(n5633), .A1(n5626), .S(n4208), .Z(n5642) );
  CMXI2X1 U14834 ( .A0(n5642), .A1(n5627), .S(n3190), .Z(n5657) );
  CMXI2X1 U14835 ( .A0(n5657), .A1(n5628), .S(n4217), .Z(n5677) );
  CMXI2X1 U14836 ( .A0(n5677), .A1(n5629), .S(n4226), .Z(n5706) );
  CMXI2X1 U14837 ( .A0(n5706), .A1(n5630), .S(n3763), .Z(n5744) );
  CND2IX1 U14838 ( .B(n5810), .A(n3730), .Z(n5912) );
  CMXI2X1 U14839 ( .A0(n5912), .A1(n5631), .S(n3845), .Z(N526) );
  CMXI2X1 U14840 ( .A0(n5641), .A1(n5633), .S(n4207), .Z(n5649) );
  CMXI2X1 U14841 ( .A0(n5649), .A1(n5634), .S(n3194), .Z(n5662) );
  CMXI2X1 U14842 ( .A0(n5662), .A1(n5635), .S(n4215), .Z(n5681) );
  CMXI2X1 U14843 ( .A0(n5681), .A1(n5636), .S(n4223), .Z(n5709) );
  CMXI2X1 U14844 ( .A0(n5709), .A1(n5637), .S(n3765), .Z(n5746) );
  CND2IX1 U14845 ( .B(n5812), .A(n3726), .Z(n5914) );
  CMXI2X1 U14846 ( .A0(n5914), .A1(n5638), .S(n3846), .Z(N527) );
  CMXI2X1 U14847 ( .A0(n5648), .A1(n5641), .S(n4208), .Z(n5656) );
  CMXI2X1 U14848 ( .A0(n5656), .A1(n5642), .S(n3192), .Z(n5667) );
  CMXI2X1 U14849 ( .A0(n5667), .A1(n5643), .S(n4219), .Z(n5685) );
  CMXI2X1 U14850 ( .A0(n5685), .A1(n5644), .S(n4222), .Z(n5712) );
  CMXI2X1 U14851 ( .A0(n5712), .A1(n5645), .S(n3762), .Z(n5748) );
  CND2IX1 U14852 ( .B(n5814), .A(n3724), .Z(n5916) );
  CMXI2X1 U14853 ( .A0(n5916), .A1(n5646), .S(n3847), .Z(N528) );
  CMXI2X1 U14854 ( .A0(n5655), .A1(n5648), .S(n4207), .Z(n5661) );
  CMXI2X1 U14855 ( .A0(n5661), .A1(n5649), .S(n3194), .Z(n5672) );
  CMXI2X1 U14856 ( .A0(n5672), .A1(n5650), .S(n4220), .Z(n5689) );
  CMXI2X1 U14857 ( .A0(n5689), .A1(n5651), .S(n4226), .Z(n5715) );
  CMXI2X1 U14858 ( .A0(n5715), .A1(n5652), .S(n3765), .Z(n5750) );
  CND2IX1 U14859 ( .B(n5816), .A(n3726), .Z(n5918) );
  CMXI2X1 U14860 ( .A0(n5918), .A1(n5653), .S(n3848), .Z(N529) );
  CMXI2X1 U14861 ( .A0(n5660), .A1(n5655), .S(n4209), .Z(n5666) );
  CMXI2X1 U14862 ( .A0(n5666), .A1(n5656), .S(n3190), .Z(n5676) );
  CMXI2X1 U14863 ( .A0(n5676), .A1(n5657), .S(n4218), .Z(n5693) );
  CMXI2X1 U14864 ( .A0(n5693), .A1(n5658), .S(n4222), .Z(n5717) );
  CMXI2X1 U14865 ( .A0(n5717), .A1(n5659), .S(n3762), .Z(n5751) );
  CMXI2X1 U14866 ( .A0(n5671), .A1(n5661), .S(n3192), .Z(n5680) );
  CMXI2X1 U14867 ( .A0(n5680), .A1(n5662), .S(n4218), .Z(n5696) );
  CMXI2X1 U14868 ( .A0(n5696), .A1(n5663), .S(n4221), .Z(n5719) );
  CMXI2X1 U14869 ( .A0(n5719), .A1(n5664), .S(n3764), .Z(n5752) );
  CMX2X1 U14870 ( .A0(n5665), .A1(n5752), .S(n3205), .Z(n5818) );
  CMXI2X1 U14871 ( .A0(n5684), .A1(n5667), .S(n4214), .Z(n5699) );
  CMXI2X1 U14872 ( .A0(n5699), .A1(n5668), .S(n4225), .Z(n5722) );
  CMXI2X1 U14873 ( .A0(n5722), .A1(n5669), .S(n3763), .Z(n5754) );
  CMX2X1 U14874 ( .A0(n5670), .A1(n5754), .S(n3205), .Z(n5819) );
  CMXI2X1 U14875 ( .A0(n5688), .A1(n5672), .S(n4217), .Z(n5702) );
  CMXI2X1 U14876 ( .A0(n5702), .A1(n5673), .S(n4226), .Z(n5724) );
  CMXI2X1 U14877 ( .A0(n5724), .A1(n5674), .S(n3766), .Z(n5756) );
  CMX2X1 U14878 ( .A0(n5675), .A1(n5756), .S(n3211), .Z(n5820) );
  CMXI2X1 U14879 ( .A0(n5705), .A1(n5677), .S(n4226), .Z(n5726) );
  CMXI2X1 U14880 ( .A0(n5726), .A1(n5678), .S(n3765), .Z(n5758) );
  CMX2X1 U14881 ( .A0(n5679), .A1(n5758), .S(n3215), .Z(n5822) );
  CMXI2X1 U14882 ( .A0(n5708), .A1(n5681), .S(n4226), .Z(n5728) );
  CMXI2X1 U14883 ( .A0(n5728), .A1(n5682), .S(n3763), .Z(n5760) );
  CMX2X1 U14884 ( .A0(n5683), .A1(n5760), .S(n3211), .Z(n5823) );
  CMXI2X1 U14885 ( .A0(n5711), .A1(n5685), .S(n4226), .Z(n5730) );
  CMXI2X1 U14886 ( .A0(n5730), .A1(n5686), .S(n3762), .Z(n5763) );
  CMX2X1 U14887 ( .A0(n5687), .A1(n5763), .S(n3209), .Z(n5824) );
  CMXI2X1 U14888 ( .A0(n5714), .A1(n5689), .S(n4226), .Z(n5732) );
  CMXI2X1 U14889 ( .A0(n5732), .A1(n5690), .S(n3763), .Z(n5765) );
  CMX2X1 U14890 ( .A0(n5691), .A1(n5765), .S(n3209), .Z(n5825) );
  CMXI2X1 U14891 ( .A0(n5734), .A1(n5694), .S(n3765), .Z(n5767) );
  CMX2X1 U14892 ( .A0(n5695), .A1(n5767), .S(n3203), .Z(n5826) );
  CMXI2X1 U14893 ( .A0(n5736), .A1(n5697), .S(n3764), .Z(n5769) );
  CMX2X1 U14894 ( .A0(n5698), .A1(n5769), .S(n3205), .Z(n5827) );
  CMXI2X1 U14895 ( .A0(n5738), .A1(n5700), .S(n3762), .Z(n5771) );
  CMX2X1 U14896 ( .A0(n5701), .A1(n5771), .S(n3201), .Z(n5828) );
  CMXI2X1 U14897 ( .A0(n5740), .A1(n5703), .S(n3766), .Z(n5773) );
  CMX2X1 U14898 ( .A0(n5704), .A1(n5773), .S(n3201), .Z(n5829) );
  CMXI2X1 U14899 ( .A0(n5743), .A1(n5706), .S(n3762), .Z(n5775) );
  CMX2X1 U14900 ( .A0(n5707), .A1(n5775), .S(n3205), .Z(n5830) );
  CMXI2X1 U14901 ( .A0(n5745), .A1(n5709), .S(n3764), .Z(n5777) );
  CMX2X1 U14902 ( .A0(n5710), .A1(n5777), .S(n3201), .Z(n5831) );
  CMXI2X1 U14903 ( .A0(n5747), .A1(n5712), .S(n3763), .Z(n5779) );
  CMX2X1 U14904 ( .A0(n5713), .A1(n5779), .S(n3213), .Z(n5833) );
  CMXI2X1 U14905 ( .A0(n5749), .A1(n5715), .S(n3764), .Z(n5781) );
  CMX2X1 U14906 ( .A0(n5716), .A1(n5781), .S(n3213), .Z(n5834) );
  CMX2X1 U14907 ( .A0(n5718), .A1(n5784), .S(n3205), .Z(n5835) );
  CMX2X1 U14908 ( .A0(n5720), .A1(n5786), .S(n3201), .Z(n5836) );
  CMX2X1 U14909 ( .A0(n5723), .A1(n5788), .S(n3215), .Z(n5837) );
  CMX2X1 U14910 ( .A0(n5725), .A1(n5790), .S(n3203), .Z(n5838) );
  CMX2X1 U14911 ( .A0(n5727), .A1(n5792), .S(n3207), .Z(n5839) );
  CMX2X1 U14912 ( .A0(n5729), .A1(n5794), .S(n3211), .Z(n5840) );
  CMX2X1 U14913 ( .A0(n5731), .A1(n5796), .S(n3201), .Z(n5841) );
  CMX2X1 U14914 ( .A0(n5733), .A1(n5798), .S(n3213), .Z(n5842) );
  CMX2X1 U14915 ( .A0(n5735), .A1(n5800), .S(n3213), .Z(n5845) );
  CMX2X1 U14916 ( .A0(n5737), .A1(n5802), .S(n3213), .Z(n5846) );
  CMX2X1 U14917 ( .A0(n5739), .A1(n5805), .S(n3215), .Z(n5847) );
  CMX2X1 U14918 ( .A0(n5741), .A1(n5807), .S(n3203), .Z(n5848) );
  CMX2X1 U14919 ( .A0(n5744), .A1(n5809), .S(n3207), .Z(n5849) );
  CMX2X1 U14920 ( .A0(n5746), .A1(n5811), .S(n3201), .Z(n5850) );
  CMX2X1 U14921 ( .A0(n5748), .A1(n5813), .S(n3199), .Z(n5851) );
  CMX2X1 U14922 ( .A0(n5750), .A1(n5815), .S(n3209), .Z(n5852) );
  CMX2X1 U14923 ( .A0(n5753), .A1(n5854), .S(n3728), .Z(n5956) );
  CMX2X1 U14924 ( .A0(n5755), .A1(n5857), .S(n3723), .Z(n5957) );
  CMX2X1 U14925 ( .A0(n5757), .A1(n5859), .S(n3723), .Z(n5958) );
  CMX2X1 U14926 ( .A0(n5759), .A1(n5861), .S(n3723), .Z(n5959) );
  CMX2X1 U14927 ( .A0(n5761), .A1(n5863), .S(n3722), .Z(n5960) );
  CMX2X1 U14928 ( .A0(n5764), .A1(n5865), .S(n3725), .Z(n5961) );
  CMX2X1 U14929 ( .A0(n5766), .A1(n5867), .S(n3725), .Z(n5962) );
  CMX2X1 U14930 ( .A0(n5768), .A1(n5869), .S(n3730), .Z(n5964) );
  CMX2X1 U14931 ( .A0(n5770), .A1(n5871), .S(n3729), .Z(n5965) );
  CMX2X1 U14932 ( .A0(n5772), .A1(n5873), .S(n3722), .Z(n5966) );
  CMX2X1 U14933 ( .A0(n5774), .A1(n5875), .S(n3724), .Z(n5967) );
  CMX2X1 U14934 ( .A0(n5776), .A1(n5878), .S(n3726), .Z(n5968) );
  CMX2X1 U14935 ( .A0(n5778), .A1(n5880), .S(n3727), .Z(n5969) );
  CMX2X1 U14936 ( .A0(n5780), .A1(n5882), .S(n3729), .Z(n5970) );
  CMX2X1 U14937 ( .A0(n5782), .A1(n5884), .S(n3724), .Z(n5971) );
  CMX2X1 U14938 ( .A0(n5785), .A1(n5886), .S(n3725), .Z(n5972) );
  CMX2X1 U14939 ( .A0(n5787), .A1(n5888), .S(n3729), .Z(n5973) );
  CMX2X1 U14940 ( .A0(n5789), .A1(n5890), .S(n3730), .Z(n5975) );
  CMX2X1 U14941 ( .A0(n5791), .A1(n5892), .S(n3729), .Z(n5976) );
  CMX2X1 U14942 ( .A0(n5793), .A1(n5894), .S(n3723), .Z(n5977) );
  CMX2X1 U14943 ( .A0(n5795), .A1(n5896), .S(n3728), .Z(n5978) );
  CMX2X1 U14944 ( .A0(n5797), .A1(n5899), .S(n3726), .Z(n5979) );
  CMX2X1 U14945 ( .A0(n5799), .A1(n5901), .S(n3724), .Z(n5980) );
  CMX2X1 U14946 ( .A0(n5801), .A1(n5903), .S(n3722), .Z(n5981) );
  CMX2X1 U14947 ( .A0(n5803), .A1(n5905), .S(n3728), .Z(n5982) );
  CMX2X1 U14948 ( .A0(n5806), .A1(n5907), .S(n3722), .Z(n5983) );
  CMX2X1 U14949 ( .A0(n5808), .A1(n5909), .S(n3724), .Z(n5984) );
  CMX2X1 U14950 ( .A0(n5810), .A1(n5911), .S(n3724), .Z(n5987) );
  CMX2X1 U14951 ( .A0(n5812), .A1(n5913), .S(n3723), .Z(n5988) );
  CMX2X1 U14952 ( .A0(n5814), .A1(n5915), .S(n3725), .Z(n5989) );
  CMX2X1 U14953 ( .A0(n5816), .A1(n5917), .S(n3727), .Z(n5990) );
  CND2IX1 U14954 ( .B(n5854), .A(n3734), .Z(n6028) );
  CMXI2X1 U14955 ( .A0(n6028), .A1(n5855), .S(n3840), .Z(N627) );
  CND2IX1 U14956 ( .B(n5857), .A(n3735), .Z(n6031) );
  CMXI2X1 U14957 ( .A0(n6031), .A1(n5858), .S(n3849), .Z(N628) );
  CND2IX1 U14958 ( .B(n5859), .A(n3735), .Z(n6035) );
  CMXI2X1 U14959 ( .A0(n6035), .A1(n5860), .S(n3850), .Z(N629) );
  CND2IX1 U14960 ( .B(n5861), .A(n3736), .Z(n6040) );
  CMXI2X1 U14961 ( .A0(n6040), .A1(n5862), .S(n3851), .Z(N630) );
  CND2IX1 U14962 ( .B(n5863), .A(n3739), .Z(n6045) );
  CMXI2X1 U14963 ( .A0(n6045), .A1(n5864), .S(n3852), .Z(N631) );
  CMXI2X1 U14964 ( .A0(n6050), .A1(n5866), .S(n3853), .Z(N632) );
  CND2IX1 U14965 ( .B(n5867), .A(n3740), .Z(n6055) );
  CMXI2X1 U14966 ( .A0(n6055), .A1(n5868), .S(n3834), .Z(N633) );
  CND2IX1 U14967 ( .B(n5869), .A(n3736), .Z(n6060) );
  CMXI2X1 U14968 ( .A0(n6060), .A1(n5870), .S(n3835), .Z(N634) );
  CND2IX1 U14969 ( .B(n5871), .A(n3733), .Z(n6066) );
  CMXI2X1 U14970 ( .A0(n6066), .A1(n5872), .S(n3836), .Z(N635) );
  CMXI2X1 U14971 ( .A0(n6071), .A1(n5874), .S(n3837), .Z(N636) );
  CND2IX1 U14972 ( .B(n5875), .A(n3731), .Z(n6076) );
  CMXI2X1 U14973 ( .A0(n6076), .A1(n5876), .S(n3838), .Z(N637) );
  CMXI2X1 U14974 ( .A0(n6080), .A1(n5879), .S(n3849), .Z(N638) );
  CND2IX1 U14975 ( .B(n5880), .A(n3738), .Z(n6084) );
  CMXI2X1 U14976 ( .A0(n6084), .A1(n5881), .S(n3841), .Z(N639) );
  CND2IX1 U14977 ( .B(n5882), .A(n3732), .Z(n6089) );
  CMXI2X1 U14978 ( .A0(n6089), .A1(n5883), .S(n3842), .Z(N640) );
  CND2IX1 U14979 ( .B(n5884), .A(n3731), .Z(n6093) );
  CMXI2X1 U14980 ( .A0(n6093), .A1(n5885), .S(n3839), .Z(N641) );
  CMXI2X1 U14981 ( .A0(n6096), .A1(n5887), .S(n3843), .Z(N642) );
  CMXI2X1 U14982 ( .A0(n6100), .A1(n5889), .S(n3839), .Z(N643) );
  CND2IX1 U14983 ( .B(n5890), .A(n3731), .Z(n6104) );
  CMXI2X1 U14984 ( .A0(n6104), .A1(n5891), .S(n3840), .Z(N644) );
  CMXI2X1 U14985 ( .A0(n6108), .A1(n5893), .S(n3841), .Z(N645) );
  CND2IX1 U14986 ( .B(n5894), .A(n3739), .Z(n6112) );
  CMXI2X1 U14987 ( .A0(n6112), .A1(n5895), .S(n3842), .Z(N646) );
  CMXI2X1 U14988 ( .A0(n6116), .A1(n5897), .S(n3841), .Z(N647) );
  CMXI2X1 U14989 ( .A0(n6120), .A1(n5900), .S(n3843), .Z(N648) );
  CMXI2X1 U14990 ( .A0(n6124), .A1(n5902), .S(n3844), .Z(N649) );
  CMXI2X1 U14991 ( .A0(n6128), .A1(n5904), .S(n3845), .Z(N650) );
  CMXI2X1 U14992 ( .A0(n6131), .A1(n5906), .S(n3846), .Z(N651) );
  CMXI2X1 U14993 ( .A0(n6134), .A1(n5908), .S(n3847), .Z(N652) );
  CMXI2X1 U14994 ( .A0(n6137), .A1(n5910), .S(n3848), .Z(N653) );
  CND2IX1 U14995 ( .B(n5911), .A(n3738), .Z(n6140) );
  CMXI2X1 U14996 ( .A0(n6140), .A1(n5912), .S(n3849), .Z(N654) );
  CMXI2X1 U14997 ( .A0(n6143), .A1(n5914), .S(n3850), .Z(N655) );
  CND2IX1 U14998 ( .B(n5915), .A(n3733), .Z(n6146) );
  CMXI2X1 U14999 ( .A0(n6146), .A1(n5916), .S(n3851), .Z(N656) );
  CMXI2X1 U15000 ( .A0(n6149), .A1(n5918), .S(n3852), .Z(N657) );
  CND2IX1 U15001 ( .B(n6228), .A(n3725), .Z(n6329) );
  CMXI2X1 U15002 ( .A0(n6329), .A1(n6028), .S(n3850), .Z(N755) );
  CMXI2X1 U15003 ( .A0(n6033), .A1(n6030), .S(n4211), .Z(n6039) );
  CND2IX1 U15004 ( .B(n6230), .A(n3722), .Z(n6331) );
  CMXI2X1 U15005 ( .A0(n6331), .A1(n6031), .S(n3844), .Z(N756) );
  CMXI2X1 U15006 ( .A0(n6038), .A1(n6033), .S(n4207), .Z(n6043) );
  CMXI2X1 U15007 ( .A0(n6043), .A1(n6034), .S(n3194), .Z(n6054) );
  CND2IX1 U15008 ( .B(n6232), .A(n3730), .Z(n6333) );
  CMXI2X1 U15009 ( .A0(n6333), .A1(n6035), .S(n3845), .Z(N757) );
  CMXI2X1 U15010 ( .A0(n6042), .A1(n6038), .S(n4210), .Z(n6048) );
  CMXI2X1 U15011 ( .A0(n6048), .A1(n6039), .S(n3188), .Z(n6059) );
  CND2IX1 U15012 ( .B(n6234), .A(n3722), .Z(n6335) );
  CMXI2X1 U15013 ( .A0(n6335), .A1(n6040), .S(n3840), .Z(N758) );
  CMXI2X1 U15014 ( .A0(n6047), .A1(n6042), .S(n4204), .Z(n6053) );
  CMXI2X1 U15015 ( .A0(n6053), .A1(n6043), .S(n3194), .Z(n6064) );
  CMXI2X1 U15016 ( .A0(n6064), .A1(n6044), .S(n4220), .Z(n6083) );
  CND2IX1 U15017 ( .B(n6236), .A(n3727), .Z(n6337) );
  CMXI2X1 U15018 ( .A0(n6337), .A1(n6045), .S(n3846), .Z(N759) );
  CMXI2X1 U15019 ( .A0(n6052), .A1(n6047), .S(n4205), .Z(n6058) );
  CMXI2X1 U15020 ( .A0(n6058), .A1(n6048), .S(n3190), .Z(n6069) );
  CMXI2X1 U15021 ( .A0(n6069), .A1(n6049), .S(n3246), .Z(n6088) );
  CMXI2X1 U15022 ( .A0(n6340), .A1(n6050), .S(n3853), .Z(N760) );
  CMXI2X1 U15023 ( .A0(n6057), .A1(n6052), .S(n4206), .Z(n6063) );
  CMXI2X1 U15024 ( .A0(n6063), .A1(n6053), .S(n3188), .Z(n6074) );
  CMXI2X1 U15025 ( .A0(n6074), .A1(n6054), .S(n3247), .Z(n6092) );
  CMXI2X1 U15026 ( .A0(n6342), .A1(n6055), .S(n3834), .Z(N761) );
  CMXI2X1 U15027 ( .A0(n6061), .A1(n6057), .S(n4209), .Z(n6067) );
  CMXI2X1 U15028 ( .A0(n6067), .A1(n6058), .S(n3192), .Z(n6077) );
  CMXI2X1 U15029 ( .A0(n6077), .A1(n6059), .S(n4219), .Z(n6094) );
  CMXI2X1 U15030 ( .A0(n6343), .A1(n6060), .S(n3835), .Z(N762) );
  CMXI2X1 U15031 ( .A0(n6062), .A1(n6061), .S(n4203), .Z(n6072) );
  CMXI2X1 U15032 ( .A0(n6072), .A1(n6063), .S(n3194), .Z(n6081) );
  CMXI2X1 U15033 ( .A0(n6081), .A1(n6064), .S(n4213), .Z(n6097) );
  CMXI2X1 U15034 ( .A0(n6097), .A1(n6065), .S(n4226), .Z(n6129) );
  CMXI2X1 U15035 ( .A0(n6345), .A1(n6066), .S(n3836), .Z(N763) );
  CMXI2X1 U15036 ( .A0(n6068), .A1(n6067), .S(n3192), .Z(n6086) );
  CMXI2X1 U15037 ( .A0(n6086), .A1(n6069), .S(n4217), .Z(n6101) );
  CMXI2X1 U15038 ( .A0(n6101), .A1(n6070), .S(n4226), .Z(n6132) );
  CMXI2X1 U15039 ( .A0(n6347), .A1(n6071), .S(n3842), .Z(N764) );
  CMXI2X1 U15040 ( .A0(n6073), .A1(n6072), .S(n3192), .Z(n6090) );
  CMXI2X1 U15041 ( .A0(n6090), .A1(n6074), .S(n4216), .Z(n6105) );
  CMXI2X1 U15042 ( .A0(n6105), .A1(n6075), .S(n4226), .Z(n6135) );
  CMXI2X1 U15043 ( .A0(n6349), .A1(n6076), .S(n3837), .Z(N765) );
  CMXI2X1 U15044 ( .A0(n6078), .A1(n6077), .S(n4219), .Z(n6109) );
  CMXI2X1 U15045 ( .A0(n6109), .A1(n6079), .S(n4226), .Z(n6138) );
  CMXI2X1 U15046 ( .A0(n6351), .A1(n6080), .S(n3838), .Z(N766) );
  CMXI2X1 U15047 ( .A0(n6082), .A1(n6081), .S(n4218), .Z(n6113) );
  CMXI2X1 U15048 ( .A0(n6113), .A1(n6083), .S(n4226), .Z(n6141) );
  CMXI2X1 U15049 ( .A0(n6353), .A1(n6084), .S(n3839), .Z(N767) );
  CMXI2X1 U15050 ( .A0(n6087), .A1(n6086), .S(n4220), .Z(n6117) );
  CMXI2X1 U15051 ( .A0(n6117), .A1(n6088), .S(n4226), .Z(n6144) );
  CMXI2X1 U15052 ( .A0(n6355), .A1(n6089), .S(n3840), .Z(N768) );
  CMXI2X1 U15053 ( .A0(n6091), .A1(n6090), .S(n4217), .Z(n6121) );
  CMXI2X1 U15054 ( .A0(n6121), .A1(n6092), .S(n4226), .Z(n6147) );
  CMXI2X1 U15055 ( .A0(n6357), .A1(n6093), .S(n3841), .Z(N769) );
  CMXI2X1 U15056 ( .A0(n6095), .A1(n6094), .S(n4225), .Z(n6150) );
  CMXI2X1 U15057 ( .A0(n6360), .A1(n6096), .S(n3842), .Z(N770) );
  CMXI2X1 U15058 ( .A0(n6098), .A1(n6097), .S(n4225), .Z(n6152) );
  CMXI2X1 U15059 ( .A0(n6152), .A1(n6099), .S(n3762), .Z(n6194) );
  CMXI2X1 U15060 ( .A0(n6362), .A1(n6100), .S(n3843), .Z(N771) );
  CMXI2X1 U15061 ( .A0(n6102), .A1(n6101), .S(n4225), .Z(n6156) );
  CMXI2X1 U15062 ( .A0(n6156), .A1(n6103), .S(n3763), .Z(n6196) );
  CMXI2X1 U15063 ( .A0(n6364), .A1(n6104), .S(n3844), .Z(N772) );
  CMXI2X1 U15064 ( .A0(n6106), .A1(n6105), .S(n4225), .Z(n6159) );
  CMXI2X1 U15065 ( .A0(n6159), .A1(n6107), .S(n3764), .Z(n6198) );
  CMXI2X1 U15066 ( .A0(n6366), .A1(n6108), .S(n3845), .Z(N773) );
  CMXI2X1 U15067 ( .A0(n6110), .A1(n6109), .S(n4224), .Z(n6162) );
  CMXI2X1 U15068 ( .A0(n6162), .A1(n6111), .S(n3762), .Z(n6200) );
  CMXI2X1 U15069 ( .A0(n6368), .A1(n6112), .S(n3846), .Z(N774) );
  CMXI2X1 U15070 ( .A0(n6114), .A1(n6113), .S(n4223), .Z(n6165) );
  CMXI2X1 U15071 ( .A0(n6165), .A1(n6115), .S(n3764), .Z(n6202) );
  CMXI2X1 U15072 ( .A0(n6370), .A1(n6116), .S(n3851), .Z(N775) );
  CMXI2X1 U15073 ( .A0(n6118), .A1(n6117), .S(n4222), .Z(n6168) );
  CMXI2X1 U15074 ( .A0(n6168), .A1(n6119), .S(n3766), .Z(n6205) );
  CMXI2X1 U15075 ( .A0(n6372), .A1(n6120), .S(n3847), .Z(N776) );
  CMXI2X1 U15076 ( .A0(n6122), .A1(n6121), .S(n4221), .Z(n6171) );
  CMXI2X1 U15077 ( .A0(n6171), .A1(n6123), .S(n3762), .Z(n6207) );
  CMXI2X1 U15078 ( .A0(n6374), .A1(n6124), .S(n3848), .Z(N777) );
  CMXI2X1 U15079 ( .A0(n6127), .A1(n6126), .S(n3766), .Z(n6209) );
  CMXI2X1 U15080 ( .A0(n6376), .A1(n6128), .S(n3841), .Z(N778) );
  CMXI2X1 U15081 ( .A0(n6130), .A1(n6129), .S(n3764), .Z(n6211) );
  CMXI2X1 U15082 ( .A0(n6378), .A1(n6131), .S(n3849), .Z(N779) );
  CMXI2X1 U15083 ( .A0(n6133), .A1(n6132), .S(n3766), .Z(n6213) );
  CMXI2X1 U15084 ( .A0(n6381), .A1(n6134), .S(n3847), .Z(N780) );
  CMXI2X1 U15085 ( .A0(n6136), .A1(n6135), .S(n3763), .Z(n6215) );
  CMXI2X1 U15086 ( .A0(n6383), .A1(n6137), .S(n3848), .Z(N781) );
  CMXI2X1 U15087 ( .A0(n6139), .A1(n6138), .S(n3764), .Z(n6217) );
  CMXI2X1 U15088 ( .A0(n6385), .A1(n6140), .S(n3849), .Z(N782) );
  CMXI2X1 U15089 ( .A0(n6142), .A1(n6141), .S(n3765), .Z(n6219) );
  CMXI2X1 U15090 ( .A0(n6387), .A1(n6143), .S(n3850), .Z(N783) );
  CMXI2X1 U15091 ( .A0(n6145), .A1(n6144), .S(n3763), .Z(n6221) );
  CMXI2X1 U15092 ( .A0(n6389), .A1(n6146), .S(n3843), .Z(N784) );
  CMXI2X1 U15093 ( .A0(n6148), .A1(n6147), .S(n3765), .Z(n6223) );
  CMXI2X1 U15094 ( .A0(n6391), .A1(n6149), .S(n3851), .Z(N785) );
  CMXI2X1 U15095 ( .A0(n6151), .A1(n6150), .S(n3766), .Z(n6226) );
  CMXI2X1 U15096 ( .A0(n6153), .A1(n6152), .S(n3765), .Z(n6227) );
  CMX2X1 U15097 ( .A0(n6154), .A1(n6227), .S(n3215), .Z(n6293) );
  CMXI2X1 U15098 ( .A0(n6157), .A1(n6156), .S(n3766), .Z(n6229) );
  CMX2X1 U15099 ( .A0(n6158), .A1(n6229), .S(n3201), .Z(n6294) );
  CMXI2X1 U15100 ( .A0(n6160), .A1(n6159), .S(n3765), .Z(n6231) );
  CMX2X1 U15101 ( .A0(n6161), .A1(n6231), .S(n3213), .Z(n6295) );
  CMXI2X1 U15102 ( .A0(n6163), .A1(n6162), .S(n3762), .Z(n6233) );
  CMX2X1 U15103 ( .A0(n6164), .A1(n6233), .S(n3205), .Z(n6296) );
  CMXI2X1 U15104 ( .A0(n6166), .A1(n6165), .S(n3764), .Z(n6235) );
  CMX2X1 U15105 ( .A0(n6167), .A1(n6235), .S(n3199), .Z(n6297) );
  CMXI2X1 U15106 ( .A0(n6169), .A1(n6168), .S(n3763), .Z(n6237) );
  CMX2X1 U15107 ( .A0(n6170), .A1(n6237), .S(n3209), .Z(n6298) );
  CMXI2X1 U15108 ( .A0(n6172), .A1(n6171), .S(n3762), .Z(n6239) );
  CMX2X1 U15109 ( .A0(n6173), .A1(n6239), .S(n3199), .Z(n6299) );
  CMX2X1 U15110 ( .A0(n6175), .A1(n6174), .S(n3205), .Z(n6301) );
  CMX2X1 U15111 ( .A0(n6177), .A1(n6176), .S(n3213), .Z(n6302) );
  CMX2X1 U15112 ( .A0(n6179), .A1(n6178), .S(n3203), .Z(n6303) );
  CMX2X1 U15113 ( .A0(n6181), .A1(n6180), .S(n3213), .Z(n6304) );
  CMX2X1 U15114 ( .A0(n6184), .A1(n6183), .S(n3199), .Z(n6305) );
  CMX2X1 U15115 ( .A0(n6186), .A1(n6185), .S(n3209), .Z(n6306) );
  CMX2X1 U15116 ( .A0(n6188), .A1(n6187), .S(n3209), .Z(n6307) );
  CMX2X1 U15117 ( .A0(n6190), .A1(n6189), .S(n3209), .Z(n6308) );
  CMX2X1 U15118 ( .A0(n6192), .A1(n6191), .S(n3211), .Z(n6309) );
  CMX2X1 U15119 ( .A0(n6194), .A1(n6193), .S(n3211), .Z(n6310) );
  CMX2X1 U15120 ( .A0(n6196), .A1(n6195), .S(n3203), .Z(n6312) );
  CMX2X1 U15121 ( .A0(n6198), .A1(n6197), .S(n3207), .Z(n6313) );
  CMX2X1 U15122 ( .A0(n6200), .A1(n6199), .S(n3215), .Z(n6314) );
  CMX2X1 U15123 ( .A0(n6202), .A1(n6201), .S(n3201), .Z(n6315) );
  CMX2X1 U15124 ( .A0(n6205), .A1(n6204), .S(n3209), .Z(n6316) );
  CMX2X1 U15125 ( .A0(n6207), .A1(n6206), .S(n3203), .Z(n6317) );
  CMX2X1 U15126 ( .A0(n6209), .A1(n6208), .S(n3213), .Z(n6318) );
  CMX2X1 U15127 ( .A0(n6211), .A1(n6210), .S(n3215), .Z(n6319) );
  CMX2X1 U15128 ( .A0(n6213), .A1(n6212), .S(n3205), .Z(n6320) );
  CMX2X1 U15129 ( .A0(n6215), .A1(n6214), .S(n3209), .Z(n6321) );
  CMX2X1 U15130 ( .A0(n6217), .A1(n6216), .S(n3201), .Z(n6323) );
  CMX2X1 U15131 ( .A0(n6219), .A1(n6218), .S(n3205), .Z(n6324) );
  CMX2X1 U15132 ( .A0(n6221), .A1(n6220), .S(n3207), .Z(n6325) );
  CMX2X1 U15133 ( .A0(n6223), .A1(n6222), .S(n3207), .Z(n6326) );
  CMX2X1 U15134 ( .A0(n6228), .A1(n6328), .S(n3724), .Z(n6430) );
  CMX2X1 U15135 ( .A0(n6230), .A1(n6330), .S(n3728), .Z(n6432) );
  CMX2X1 U15136 ( .A0(n6232), .A1(n6332), .S(n3727), .Z(n6433) );
  CMX2X1 U15137 ( .A0(n6234), .A1(n6334), .S(n3724), .Z(n6434) );
  CMX2X1 U15138 ( .A0(n6236), .A1(n6336), .S(n3723), .Z(n6435) );
  CMX2X1 U15139 ( .A0(n6238), .A1(n6339), .S(n3730), .Z(n6436) );
  CMX2X1 U15140 ( .A0(n6240), .A1(n6341), .S(n3722), .Z(n6437) );
  CMXI2X1 U15141 ( .A0(n6242), .A1(n6241), .S(n3722), .Z(n6438) );
  CMXI2X1 U15142 ( .A0(n6244), .A1(n6243), .S(n3725), .Z(n6439) );
  CMXI2X1 U15143 ( .A0(n6247), .A1(n6246), .S(n3723), .Z(n6440) );
  CMXI2X1 U15144 ( .A0(n6249), .A1(n6248), .S(n3728), .Z(n6441) );
  CMXI2X1 U15145 ( .A0(n6251), .A1(n6250), .S(n3726), .Z(n6443) );
  CMXI2X1 U15146 ( .A0(n6253), .A1(n6252), .S(n3722), .Z(n6444) );
  CMXI2X1 U15147 ( .A0(n6255), .A1(n6254), .S(n3728), .Z(n6445) );
  CMXI2X1 U15148 ( .A0(n6257), .A1(n6256), .S(n3729), .Z(n6446) );
  CMXI2X1 U15149 ( .A0(n6259), .A1(n6258), .S(n3724), .Z(n6447) );
  CMXI2X1 U15150 ( .A0(n6261), .A1(n6260), .S(n3721), .Z(n6448) );
  CMXI2X1 U15151 ( .A0(n6263), .A1(n6262), .S(n3730), .Z(n6449) );
  CMXI2X1 U15152 ( .A0(n6265), .A1(n6264), .S(n3728), .Z(n6450) );
  CMXI2X1 U15153 ( .A0(n6268), .A1(n6267), .S(n3725), .Z(n6451) );
  CMXI2X1 U15154 ( .A0(n6270), .A1(n6269), .S(n3725), .Z(n6452) );
  CMXI2X1 U15155 ( .A0(n6272), .A1(n6271), .S(n3723), .Z(n6454) );
  CMXI2X1 U15156 ( .A0(n6274), .A1(n6273), .S(n3726), .Z(n6455) );
  CMXI2X1 U15157 ( .A0(n6276), .A1(n6275), .S(n3728), .Z(n6456) );
  CMXI2X1 U15158 ( .A0(n6278), .A1(n6277), .S(n3729), .Z(n6457) );
  CMXI2X1 U15159 ( .A0(n6280), .A1(n6279), .S(n3725), .Z(n6458) );
  CMXI2X1 U15160 ( .A0(n6282), .A1(n6281), .S(n3725), .Z(n6459) );
  CMXI2X1 U15161 ( .A0(n6284), .A1(n6283), .S(n3728), .Z(n6460) );
  CMXI2X1 U15162 ( .A0(n6286), .A1(n6285), .S(n3728), .Z(n6461) );
  CMXI2X1 U15163 ( .A0(n6289), .A1(n6288), .S(n3724), .Z(n6462) );
  CMXI2X1 U15164 ( .A0(n6291), .A1(n6290), .S(n3723), .Z(n6463) );
  CND2IX1 U15165 ( .B(n6328), .A(n3738), .Z(n6505) );
  CMXI2X1 U15166 ( .A0(n6505), .A1(n6329), .S(n3852), .Z(N883) );
  CND2IX1 U15167 ( .B(n6330), .A(n3731), .Z(n6506) );
  CMXI2X1 U15168 ( .A0(n6506), .A1(n6331), .S(n3853), .Z(N884) );
  CND2IX1 U15169 ( .B(n6332), .A(n3732), .Z(n6507) );
  CMXI2X1 U15170 ( .A0(n6507), .A1(n6333), .S(n3834), .Z(N885) );
  CND2IX1 U15171 ( .B(n6334), .A(n3734), .Z(n6508) );
  CMXI2X1 U15172 ( .A0(n6508), .A1(n6335), .S(n3835), .Z(N886) );
  CND2IX1 U15173 ( .B(n6336), .A(n3737), .Z(n6509) );
  CMXI2X1 U15174 ( .A0(n6509), .A1(n6337), .S(n3836), .Z(N887) );
  CND2IX1 U15175 ( .B(n6339), .A(n3735), .Z(n6510) );
  CMXI2X1 U15176 ( .A0(n6510), .A1(n6340), .S(n3837), .Z(N888) );
  CND2IX1 U15177 ( .B(n6341), .A(n3733), .Z(n6511) );
  CMXI2X1 U15178 ( .A0(n6511), .A1(n6342), .S(n3838), .Z(N889) );
  CMXI2X1 U15179 ( .A0(n6344), .A1(n6343), .S(n3839), .Z(N890) );
  CMXI2X1 U15180 ( .A0(n6346), .A1(n6345), .S(n3840), .Z(N891) );
  CMXI2X1 U15181 ( .A0(n6348), .A1(n6347), .S(n3852), .Z(N892) );
  CMXI2X1 U15182 ( .A0(n6350), .A1(n6349), .S(n3850), .Z(N893) );
  CMXI2X1 U15183 ( .A0(n6352), .A1(n6351), .S(n3851), .Z(N894) );
  CMXI2X1 U15184 ( .A0(n6354), .A1(n6353), .S(n3842), .Z(N895) );
  CMXI2X1 U15185 ( .A0(n6356), .A1(n6355), .S(n3852), .Z(N896) );
  CMXI2X1 U15186 ( .A0(n6358), .A1(n6357), .S(n3841), .Z(N897) );
  CMXI2X1 U15187 ( .A0(n6361), .A1(n6360), .S(n3842), .Z(N898) );
  CMXI2X1 U15188 ( .A0(n6363), .A1(n6362), .S(n3843), .Z(N899) );
  CMXI2X1 U15189 ( .A0(n6365), .A1(n6364), .S(n3844), .Z(N900) );
  CMXI2X1 U15190 ( .A0(n6367), .A1(n6366), .S(n3844), .Z(N901) );
  CMXI2X1 U15191 ( .A0(n6369), .A1(n6368), .S(n3845), .Z(N902) );
  CMXI2X1 U15192 ( .A0(n6371), .A1(n6370), .S(n3846), .Z(N903) );
  CMXI2X1 U15193 ( .A0(n6373), .A1(n6372), .S(n3847), .Z(N904) );
  CMXI2X1 U15194 ( .A0(n6375), .A1(n6374), .S(n3848), .Z(N905) );
  CMXI2X1 U15195 ( .A0(n6377), .A1(n6376), .S(n3849), .Z(N906) );
  CMXI2X1 U15196 ( .A0(n6379), .A1(n6378), .S(n3850), .Z(N907) );
  CMXI2X1 U15197 ( .A0(n6382), .A1(n6381), .S(n3851), .Z(N908) );
  CMXI2X1 U15198 ( .A0(n6384), .A1(n6383), .S(n3852), .Z(N909) );
  CMXI2X1 U15199 ( .A0(n6386), .A1(n6385), .S(n3853), .Z(N910) );
  CMXI2X1 U15200 ( .A0(n6388), .A1(n6387), .S(n3834), .Z(N911) );
  CMXI2X1 U15201 ( .A0(n6390), .A1(n6389), .S(n3838), .Z(N912) );
  CMXI2X1 U15202 ( .A0(n6392), .A1(n6391), .S(n3839), .Z(N913) );
  CND2IX1 U15203 ( .B(n6486), .A(n3725), .Z(n6487) );
  CMXI2X1 U15204 ( .A0(n6488), .A1(n6487), .S(n3840), .Z(N115) );
  CND2IX1 U15205 ( .B(n6499), .A(n3728), .Z(n6500) );
  CMXI2X1 U15206 ( .A0(n6501), .A1(n6500), .S(n3841), .Z(N116) );
  CND2IX1 U15207 ( .B(n6512), .A(n3729), .Z(n6513) );
  CMXI2X1 U15208 ( .A0(n6514), .A1(n6513), .S(n3842), .Z(N117) );
  CMXI2X1 U15209 ( .A0(mem_data1[7]), .A1(mem_data1[6]), .S(n3890), .Z(n7256)
         );
  CMXI2X1 U15210 ( .A0(mem_data1[5]), .A1(mem_data1[4]), .S(n3890), .Z(n7259)
         );
  CMXI2X1 U15211 ( .A0(n7256), .A1(n7259), .S(n4074), .Z(n7931) );
  CMXI2X1 U15212 ( .A0(mem_data1[2]), .A1(mem_data1[3]), .S(n3866), .Z(n7258)
         );
  CMXI2X1 U15213 ( .A0(mem_data1[1]), .A1(mem_data1[0]), .S(n3888), .Z(n6516)
         );
  CMXI2X1 U15214 ( .A0(n7258), .A1(n6516), .S(n4074), .Z(n6517) );
  CMXI2X1 U15215 ( .A0(n7931), .A1(n6517), .S(n3782), .Z(n6518) );
  CMX2X1 U15216 ( .A0(mem_data1[10]), .A1(mem_data1[11]), .S(n3875), .Z(n6613)
         );
  CMXI2X1 U15217 ( .A0(mem_data1[9]), .A1(mem_data1[8]), .S(n3885), .Z(n7257)
         );
  CMXI2X1 U15218 ( .A0(n6613), .A1(n4429), .S(n4074), .Z(n7930) );
  CMX2X1 U15219 ( .A0(mem_data1[14]), .A1(mem_data1[15]), .S(n3878), .Z(n6615)
         );
  CMX2X1 U15220 ( .A0(mem_data1[12]), .A1(mem_data1[13]), .S(n3876), .Z(n6614)
         );
  CMXI2X1 U15221 ( .A0(n6615), .A1(n6614), .S(n4074), .Z(n6678) );
  CMX2X1 U15222 ( .A0(n7930), .A1(n6678), .S(n4368), .Z(n9269) );
  CMXI2X1 U15223 ( .A0(n6518), .A1(n9269), .S(n3499), .Z(N2076) );
  CMX2X1 U15224 ( .A0(mem_data1[1002]), .A1(mem_data1[1003]), .S(n3879), .Z(
        n6519) );
  CMX2X1 U15225 ( .A0(mem_data1[1000]), .A1(mem_data1[1001]), .S(n3878), .Z(
        n9547) );
  CMXI2X1 U15226 ( .A0(n6519), .A1(n9547), .S(n4074), .Z(n9554) );
  CMX2X1 U15227 ( .A0(mem_data1[1006]), .A1(mem_data1[1007]), .S(n3879), .Z(
        n6521) );
  CMX2X1 U15228 ( .A0(mem_data1[1004]), .A1(mem_data1[1005]), .S(n3880), .Z(
        n6520) );
  CMXI2X1 U15229 ( .A0(n6521), .A1(n6520), .S(n4074), .Z(n6534) );
  CMX2X1 U15230 ( .A0(n9554), .A1(n6534), .S(n4368), .Z(n9568) );
  CMX2X1 U15231 ( .A0(mem_data1[1010]), .A1(mem_data1[1011]), .S(n3881), .Z(
        n6523) );
  CMX2X1 U15232 ( .A0(mem_data1[1008]), .A1(mem_data1[1009]), .S(n3876), .Z(
        n6522) );
  CMXI2X1 U15233 ( .A0(n6523), .A1(n6522), .S(n4073), .Z(n6533) );
  CMX2X1 U15234 ( .A0(mem_data1[1014]), .A1(mem_data1[1015]), .S(n3877), .Z(
        n6525) );
  CMX2X1 U15235 ( .A0(mem_data1[1012]), .A1(mem_data1[1013]), .S(n3878), .Z(
        n6524) );
  CMXI2X1 U15236 ( .A0(n6525), .A1(n6524), .S(n4073), .Z(n6536) );
  CMX2X1 U15237 ( .A0(n6533), .A1(n6536), .S(n4368), .Z(n6551) );
  CMXI2X1 U15238 ( .A0(n9568), .A1(n6551), .S(n3465), .Z(N3076) );
  CMX2X1 U15239 ( .A0(mem_data1[1003]), .A1(mem_data1[1004]), .S(n3879), .Z(
        n6526) );
  CMX2X1 U15240 ( .A0(mem_data1[1001]), .A1(mem_data1[1002]), .S(n3869), .Z(
        n9551) );
  CMXI2X1 U15241 ( .A0(n6526), .A1(n9551), .S(n4073), .Z(n9557) );
  CMX2X1 U15242 ( .A0(mem_data1[1007]), .A1(mem_data1[1008]), .S(n3870), .Z(
        n6528) );
  CMX2X1 U15243 ( .A0(mem_data1[1005]), .A1(mem_data1[1006]), .S(n3871), .Z(
        n6527) );
  CMXI2X1 U15244 ( .A0(n6528), .A1(n6527), .S(n4073), .Z(n6538) );
  CMX2X1 U15245 ( .A0(n9557), .A1(n6538), .S(n4368), .Z(n9570) );
  CMX2X1 U15246 ( .A0(mem_data1[1011]), .A1(mem_data1[1012]), .S(n3872), .Z(
        n6530) );
  CMX2X1 U15247 ( .A0(mem_data1[1009]), .A1(mem_data1[1010]), .S(n3870), .Z(
        n6529) );
  CMXI2X1 U15248 ( .A0(n6530), .A1(n6529), .S(n4073), .Z(n6537) );
  CMX2X1 U15249 ( .A0(mem_data1[1015]), .A1(mem_data1[1016]), .S(n3862), .Z(
        n6532) );
  CMX2X1 U15250 ( .A0(mem_data1[1013]), .A1(mem_data1[1014]), .S(n3863), .Z(
        n6531) );
  CMXI2X1 U15251 ( .A0(n6532), .A1(n6531), .S(n4073), .Z(n6540) );
  CMX2X1 U15252 ( .A0(n6537), .A1(n6540), .S(n4368), .Z(n6554) );
  CMXI2X1 U15253 ( .A0(n9570), .A1(n6554), .S(n3492), .Z(N3077) );
  CMXI2X1 U15254 ( .A0(n6520), .A1(n6519), .S(n4073), .Z(n9562) );
  CMXI2X1 U15255 ( .A0(n6522), .A1(n6521), .S(n4073), .Z(n6542) );
  CMX2X1 U15256 ( .A0(n9562), .A1(n6542), .S(n4368), .Z(n9572) );
  CMXI2X1 U15257 ( .A0(n6524), .A1(n6523), .S(n4073), .Z(n6541) );
  CMX2X1 U15258 ( .A0(mem_data1[1016]), .A1(mem_data1[1017]), .S(n3862), .Z(
        n6535) );
  CMXI2X1 U15259 ( .A0(n6535), .A1(n6525), .S(n4073), .Z(n6544) );
  CMX2X1 U15260 ( .A0(n6541), .A1(n6544), .S(n4368), .Z(n6557) );
  CMXI2X1 U15261 ( .A0(n9572), .A1(n6557), .S(n3484), .Z(N3078) );
  CMXI2X1 U15262 ( .A0(n6527), .A1(n6526), .S(n4073), .Z(n9565) );
  CMXI2X1 U15263 ( .A0(n6529), .A1(n6528), .S(n4073), .Z(n6546) );
  CMX2X1 U15264 ( .A0(n9565), .A1(n6546), .S(n4368), .Z(n9574) );
  CMXI2X1 U15265 ( .A0(n6531), .A1(n6530), .S(n4073), .Z(n6545) );
  CMX2X1 U15266 ( .A0(mem_data1[1017]), .A1(mem_data1[1018]), .S(n3863), .Z(
        n6539) );
  CMXI2X1 U15267 ( .A0(n6539), .A1(n6532), .S(n4073), .Z(n6548) );
  CMX2X1 U15268 ( .A0(n6545), .A1(n6548), .S(n4368), .Z(n6560) );
  CMXI2X1 U15269 ( .A0(n9574), .A1(n6560), .S(n3484), .Z(N3079) );
  CMX2X1 U15270 ( .A0(n6534), .A1(n6533), .S(n4368), .Z(n9576) );
  CMX2X1 U15271 ( .A0(mem_data1[1018]), .A1(mem_data1[1019]), .S(n3864), .Z(
        n6543) );
  CMXI2X1 U15272 ( .A0(n6543), .A1(n6535), .S(n4073), .Z(n6550) );
  CMX2X1 U15273 ( .A0(n6536), .A1(n6550), .S(n4367), .Z(n6562) );
  CMXI2X1 U15274 ( .A0(n9576), .A1(n6562), .S(n3483), .Z(N3080) );
  CMX2X1 U15275 ( .A0(n6538), .A1(n6537), .S(n4367), .Z(n9578) );
  CMX2X1 U15276 ( .A0(mem_data1[1019]), .A1(mem_data1[1020]), .S(n3865), .Z(
        n6547) );
  CMXI2X1 U15277 ( .A0(n6547), .A1(n6539), .S(n4073), .Z(n6553) );
  CMX2X1 U15278 ( .A0(n6540), .A1(n6553), .S(n4367), .Z(n6564) );
  CMXI2X1 U15279 ( .A0(n9578), .A1(n6564), .S(n3483), .Z(N3081) );
  CMX2X1 U15280 ( .A0(n6542), .A1(n6541), .S(n4367), .Z(n9580) );
  CMX2X1 U15281 ( .A0(mem_data1[1020]), .A1(mem_data1[1021]), .S(n3880), .Z(
        n6549) );
  CMXI2X1 U15282 ( .A0(n6549), .A1(n6543), .S(n4072), .Z(n6556) );
  CMX2X1 U15283 ( .A0(n6544), .A1(n6556), .S(n4367), .Z(n6566) );
  CMXI2X1 U15284 ( .A0(n9580), .A1(n6566), .S(n3483), .Z(N3082) );
  CMX2X1 U15285 ( .A0(n6546), .A1(n6545), .S(n4367), .Z(n9582) );
  CMX2X1 U15286 ( .A0(mem_data1[1021]), .A1(mem_data1[1022]), .S(n3881), .Z(
        n6552) );
  CMXI2X1 U15287 ( .A0(n6552), .A1(n6547), .S(n4072), .Z(n6559) );
  CMX2X1 U15288 ( .A0(n6548), .A1(n6559), .S(n4367), .Z(n6568) );
  CMXI2X1 U15289 ( .A0(n9582), .A1(n6568), .S(n3483), .Z(N3083) );
  CMX2X1 U15290 ( .A0(mem_data1[1022]), .A1(mem_data1[1023]), .S(n3879), .Z(
        n6555) );
  CMXI2X1 U15291 ( .A0(n6555), .A1(n6549), .S(n4072), .Z(n6561) );
  CMX2X1 U15292 ( .A0(n6550), .A1(n6561), .S(n4367), .Z(n6569) );
  CMXI2X1 U15293 ( .A0(n6551), .A1(n6569), .S(n3483), .Z(N3084) );
  CMXI2X1 U15294 ( .A0(n6558), .A1(n6552), .S(n4072), .Z(n6563) );
  CMX2X1 U15295 ( .A0(n6553), .A1(n6563), .S(n4367), .Z(n6570) );
  CMXI2X1 U15296 ( .A0(n6554), .A1(n6570), .S(n3483), .Z(N3085) );
  CMX2X1 U15297 ( .A0(mem_data1[102]), .A1(mem_data1[103]), .S(n3864), .Z(
        n6577) );
  CMX2X1 U15298 ( .A0(mem_data1[100]), .A1(mem_data1[101]), .S(n3865), .Z(
        n9165) );
  CMXI2X1 U15299 ( .A0(n6577), .A1(n9165), .S(n4072), .Z(n9232) );
  CMX2X1 U15300 ( .A0(mem_data1[106]), .A1(mem_data1[107]), .S(n3866), .Z(
        n6579) );
  CMX2X1 U15301 ( .A0(mem_data1[104]), .A1(mem_data1[105]), .S(n3867), .Z(
        n6578) );
  CMXI2X1 U15302 ( .A0(n6579), .A1(n6578), .S(n4072), .Z(n6592) );
  CMX2X1 U15303 ( .A0(n9232), .A1(n6592), .S(n4367), .Z(n9366) );
  CMX2X1 U15304 ( .A0(mem_data1[110]), .A1(mem_data1[111]), .S(n3868), .Z(
        n6581) );
  CMX2X1 U15305 ( .A0(mem_data1[108]), .A1(mem_data1[109]), .S(n3880), .Z(
        n6580) );
  CMXI2X1 U15306 ( .A0(n6581), .A1(n6580), .S(n4072), .Z(n6591) );
  CMX2X1 U15307 ( .A0(mem_data1[114]), .A1(mem_data1[115]), .S(n3881), .Z(
        n6583) );
  CMX2X1 U15308 ( .A0(mem_data1[112]), .A1(mem_data1[113]), .S(n3869), .Z(
        n6582) );
  CMXI2X1 U15309 ( .A0(n6583), .A1(n6582), .S(n4072), .Z(n6594) );
  CMX2X1 U15310 ( .A0(n6591), .A1(n6594), .S(n4367), .Z(n6609) );
  CMXI2X1 U15311 ( .A0(n9366), .A1(n6609), .S(n3483), .Z(N2176) );
  CMX2X1 U15312 ( .A0(n6556), .A1(n6565), .S(n4366), .Z(n6571) );
  CMXI2X1 U15313 ( .A0(n6557), .A1(n6571), .S(n3483), .Z(N3086) );
  CMX2X1 U15314 ( .A0(n6559), .A1(n6567), .S(n4366), .Z(n6572) );
  CMXI2X1 U15315 ( .A0(n6560), .A1(n6572), .S(n3483), .Z(N3087) );
  CND2IX1 U15316 ( .B(n6561), .A(n3782), .Z(n6573) );
  CMXI2X1 U15317 ( .A0(n6562), .A1(n6573), .S(n3483), .Z(N3088) );
  CND2IX1 U15318 ( .B(n6563), .A(n3798), .Z(n6574) );
  CMXI2X1 U15319 ( .A0(n6564), .A1(n6574), .S(n3483), .Z(N3089) );
  CND2IX1 U15320 ( .B(n6565), .A(n3788), .Z(n6575) );
  CMXI2X1 U15321 ( .A0(n6566), .A1(n6575), .S(n3482), .Z(N3090) );
  CND2IX1 U15322 ( .B(n6567), .A(n3782), .Z(n6576) );
  CMXI2X1 U15323 ( .A0(n6568), .A1(n6576), .S(n3482), .Z(N3091) );
  CMX2X1 U15324 ( .A0(mem_data1[103]), .A1(mem_data1[104]), .S(n3870), .Z(
        n6584) );
  CMX2X1 U15325 ( .A0(mem_data1[101]), .A1(mem_data1[102]), .S(n3880), .Z(
        n9199) );
  CMXI2X1 U15326 ( .A0(n6584), .A1(n9199), .S(n4072), .Z(n9265) );
  CMX2X1 U15327 ( .A0(mem_data1[107]), .A1(mem_data1[108]), .S(n3881), .Z(
        n6586) );
  CMX2X1 U15328 ( .A0(mem_data1[105]), .A1(mem_data1[106]), .S(n3862), .Z(
        n6585) );
  CMXI2X1 U15329 ( .A0(n6586), .A1(n6585), .S(n4072), .Z(n6596) );
  CMX2X1 U15330 ( .A0(n9265), .A1(n6596), .S(n4366), .Z(n9398) );
  CMX2X1 U15331 ( .A0(mem_data1[111]), .A1(mem_data1[112]), .S(n3863), .Z(
        n6588) );
  CMX2X1 U15332 ( .A0(mem_data1[109]), .A1(mem_data1[110]), .S(n3873), .Z(
        n6587) );
  CMXI2X1 U15333 ( .A0(n6588), .A1(n6587), .S(n4072), .Z(n6595) );
  CMX2X1 U15334 ( .A0(mem_data1[115]), .A1(mem_data1[116]), .S(n3874), .Z(
        n6590) );
  CMX2X1 U15335 ( .A0(mem_data1[113]), .A1(mem_data1[114]), .S(n3875), .Z(
        n6589) );
  CMXI2X1 U15336 ( .A0(n6590), .A1(n6589), .S(n4072), .Z(n6598) );
  CMX2X1 U15337 ( .A0(n6595), .A1(n6598), .S(n4366), .Z(n6612) );
  CMXI2X1 U15338 ( .A0(n9398), .A1(n6612), .S(n3486), .Z(N2177) );
  CMXI2X1 U15339 ( .A0(n6578), .A1(n6577), .S(n4072), .Z(n9300) );
  CMXI2X1 U15340 ( .A0(n6580), .A1(n6579), .S(n4072), .Z(n6600) );
  CMX2X1 U15341 ( .A0(n9300), .A1(n6600), .S(n4366), .Z(n9430) );
  CMXI2X1 U15342 ( .A0(n6582), .A1(n6581), .S(n4072), .Z(n6599) );
  CMX2X1 U15343 ( .A0(mem_data1[116]), .A1(mem_data1[117]), .S(n3876), .Z(
        n6593) );
  CMXI2X1 U15344 ( .A0(n6593), .A1(n6583), .S(n4072), .Z(n6602) );
  CMX2X1 U15345 ( .A0(n6599), .A1(n6602), .S(n4366), .Z(n6618) );
  CMXI2X1 U15346 ( .A0(n9430), .A1(n6618), .S(n3485), .Z(N2178) );
  CMXI2X1 U15347 ( .A0(n6585), .A1(n6584), .S(n4071), .Z(n9333) );
  CMXI2X1 U15348 ( .A0(n6587), .A1(n6586), .S(n4071), .Z(n6604) );
  CMX2X1 U15349 ( .A0(n9333), .A1(n6604), .S(n4366), .Z(n9462) );
  CMXI2X1 U15350 ( .A0(n6589), .A1(n6588), .S(n4071), .Z(n6603) );
  CMX2X1 U15351 ( .A0(mem_data1[117]), .A1(mem_data1[118]), .S(n3871), .Z(
        n6597) );
  CMXI2X1 U15352 ( .A0(n6597), .A1(n6590), .S(n4071), .Z(n6606) );
  CMX2X1 U15353 ( .A0(n6603), .A1(n6606), .S(n4366), .Z(n6621) );
  CMXI2X1 U15354 ( .A0(n9462), .A1(n6621), .S(n3485), .Z(N2179) );
  CMX2X1 U15355 ( .A0(n6592), .A1(n6591), .S(n4366), .Z(n9494) );
  CMX2X1 U15356 ( .A0(mem_data1[118]), .A1(mem_data1[119]), .S(n3871), .Z(
        n6601) );
  CMXI2X1 U15357 ( .A0(n6601), .A1(n6593), .S(n4071), .Z(n6608) );
  CMX2X1 U15358 ( .A0(n6594), .A1(n6608), .S(n4366), .Z(n6624) );
  CMXI2X1 U15359 ( .A0(n9494), .A1(n6624), .S(n3485), .Z(N2180) );
  CMX2X1 U15360 ( .A0(n6596), .A1(n6595), .S(n4366), .Z(n9526) );
  CMX2X1 U15361 ( .A0(mem_data1[119]), .A1(mem_data1[120]), .S(n3872), .Z(
        n6605) );
  CMXI2X1 U15362 ( .A0(n6605), .A1(n6597), .S(n4071), .Z(n6611) );
  CMX2X1 U15363 ( .A0(n6598), .A1(n6611), .S(n4365), .Z(n6627) );
  CMXI2X1 U15364 ( .A0(n9526), .A1(n6627), .S(n3485), .Z(N2181) );
  CMX2X1 U15365 ( .A0(n6600), .A1(n6599), .S(n4365), .Z(n9560) );
  CMX2X1 U15366 ( .A0(mem_data1[120]), .A1(mem_data1[121]), .S(n3873), .Z(
        n6607) );
  CMXI2X1 U15367 ( .A0(n6607), .A1(n6601), .S(n4071), .Z(n6617) );
  CMX2X1 U15368 ( .A0(n6602), .A1(n6617), .S(n4365), .Z(n6630) );
  CMXI2X1 U15369 ( .A0(n9560), .A1(n6630), .S(n3485), .Z(N2182) );
  CMX2X1 U15370 ( .A0(n6604), .A1(n6603), .S(n4365), .Z(n9584) );
  CMX2X1 U15371 ( .A0(mem_data1[121]), .A1(mem_data1[122]), .S(n3874), .Z(
        n6610) );
  CMXI2X1 U15372 ( .A0(n6610), .A1(n6605), .S(n4071), .Z(n6620) );
  CMX2X1 U15373 ( .A0(n6606), .A1(n6620), .S(n4365), .Z(n6633) );
  CMXI2X1 U15374 ( .A0(n9584), .A1(n6633), .S(n3485), .Z(N2183) );
  CMX2X1 U15375 ( .A0(mem_data1[122]), .A1(mem_data1[123]), .S(n3875), .Z(
        n6616) );
  CMXI2X1 U15376 ( .A0(n6616), .A1(n6607), .S(n4071), .Z(n6623) );
  CMX2X1 U15377 ( .A0(n6608), .A1(n6623), .S(n4365), .Z(n6636) );
  CMXI2X1 U15378 ( .A0(n6609), .A1(n6636), .S(n3485), .Z(N2184) );
  CMX2X1 U15379 ( .A0(mem_data1[123]), .A1(mem_data1[124]), .S(n3876), .Z(
        n6619) );
  CMXI2X1 U15380 ( .A0(n6619), .A1(n6610), .S(n4071), .Z(n6626) );
  CMX2X1 U15381 ( .A0(n6611), .A1(n6626), .S(n4365), .Z(n6639) );
  CMXI2X1 U15382 ( .A0(n6612), .A1(n6639), .S(n3485), .Z(N2185) );
  CMXI2X1 U15383 ( .A0(n6614), .A1(n6613), .S(n4071), .Z(n8598) );
  CMX2X1 U15384 ( .A0(mem_data1[16]), .A1(mem_data1[17]), .S(n3877), .Z(n6676)
         );
  CMXI2X1 U15385 ( .A0(n6676), .A1(n6615), .S(n4071), .Z(n6750) );
  CMX2X1 U15386 ( .A0(n8598), .A1(n6750), .S(n4365), .Z(n7261) );
  CMX2X1 U15387 ( .A0(mem_data1[20]), .A1(mem_data1[21]), .S(n3875), .Z(n6679)
         );
  CMX2X1 U15388 ( .A0(mem_data1[18]), .A1(mem_data1[19]), .S(n3876), .Z(n6677)
         );
  CMXI2X1 U15389 ( .A0(n6679), .A1(n6677), .S(n4071), .Z(n6749) );
  CMX2X1 U15390 ( .A0(mem_data1[24]), .A1(mem_data1[25]), .S(n3877), .Z(n6681)
         );
  CMX2X1 U15391 ( .A0(mem_data1[22]), .A1(mem_data1[23]), .S(n3878), .Z(n6680)
         );
  CMXI2X1 U15392 ( .A0(n6681), .A1(n6680), .S(n4071), .Z(n6752) );
  CMX2X1 U15393 ( .A0(n6749), .A1(n6752), .S(n4365), .Z(n6887) );
  CMXI2X1 U15394 ( .A0(n7261), .A1(n6887), .S(n3485), .Z(N2086) );
  CMX2X1 U15395 ( .A0(mem_data1[124]), .A1(mem_data1[125]), .S(n3879), .Z(
        n6622) );
  CMXI2X1 U15396 ( .A0(n6622), .A1(n6616), .S(n4071), .Z(n6629) );
  CMX2X1 U15397 ( .A0(n6617), .A1(n6629), .S(n4365), .Z(n6642) );
  CMXI2X1 U15398 ( .A0(n6618), .A1(n6642), .S(n3485), .Z(N2186) );
  CMX2X1 U15399 ( .A0(mem_data1[125]), .A1(mem_data1[126]), .S(n3880), .Z(
        n6625) );
  CMXI2X1 U15400 ( .A0(n6625), .A1(n6619), .S(n4071), .Z(n6632) );
  CMX2X1 U15401 ( .A0(n6620), .A1(n6632), .S(n4365), .Z(n6645) );
  CMXI2X1 U15402 ( .A0(n6621), .A1(n6645), .S(n3485), .Z(N2187) );
  CMX2X1 U15403 ( .A0(mem_data1[126]), .A1(mem_data1[127]), .S(n3881), .Z(
        n6628) );
  CMXI2X1 U15404 ( .A0(n6628), .A1(n6622), .S(n4070), .Z(n6635) );
  CMX2X1 U15405 ( .A0(n6623), .A1(n6635), .S(n3808), .Z(n6648) );
  CMXI2X1 U15406 ( .A0(n6624), .A1(n6648), .S(n3484), .Z(N2188) );
  CMX2X1 U15407 ( .A0(mem_data1[127]), .A1(mem_data1[128]), .S(n3878), .Z(
        n6631) );
  CMXI2X1 U15408 ( .A0(n6631), .A1(n6625), .S(n4070), .Z(n6638) );
  CMX2X1 U15409 ( .A0(n6626), .A1(n6638), .S(n3809), .Z(n6651) );
  CMXI2X1 U15410 ( .A0(n6627), .A1(n6651), .S(n3484), .Z(N2189) );
  CMX2X1 U15411 ( .A0(mem_data1[128]), .A1(mem_data1[129]), .S(n3879), .Z(
        n6634) );
  CMXI2X1 U15412 ( .A0(n6634), .A1(n6628), .S(n4070), .Z(n6641) );
  CMX2X1 U15413 ( .A0(n6629), .A1(n6641), .S(n3810), .Z(n6654) );
  CMXI2X1 U15414 ( .A0(n6630), .A1(n6654), .S(n3484), .Z(N2190) );
  CMX2X1 U15415 ( .A0(mem_data1[129]), .A1(mem_data1[130]), .S(n3862), .Z(
        n6637) );
  CMXI2X1 U15416 ( .A0(n6637), .A1(n6631), .S(n4070), .Z(n6644) );
  CMX2X1 U15417 ( .A0(n6632), .A1(n6644), .S(n3811), .Z(n6657) );
  CMXI2X1 U15418 ( .A0(n6633), .A1(n6657), .S(n3484), .Z(N2191) );
  CMX2X1 U15419 ( .A0(mem_data1[130]), .A1(mem_data1[131]), .S(n3863), .Z(
        n6640) );
  CMXI2X1 U15420 ( .A0(n6640), .A1(n6634), .S(n4070), .Z(n6647) );
  CMX2X1 U15421 ( .A0(n6635), .A1(n6647), .S(n3812), .Z(n6660) );
  CMXI2X1 U15422 ( .A0(n6636), .A1(n6660), .S(n3484), .Z(N2192) );
  CMX2X1 U15423 ( .A0(mem_data1[131]), .A1(mem_data1[132]), .S(n3880), .Z(
        n6643) );
  CMXI2X1 U15424 ( .A0(n6643), .A1(n6637), .S(n4070), .Z(n6650) );
  CMX2X1 U15425 ( .A0(n6638), .A1(n6650), .S(n4357), .Z(n6663) );
  CMXI2X1 U15426 ( .A0(n6639), .A1(n6663), .S(n3484), .Z(N2193) );
  CMX2X1 U15427 ( .A0(mem_data1[132]), .A1(mem_data1[133]), .S(n3881), .Z(
        n6646) );
  CMXI2X1 U15428 ( .A0(n6646), .A1(n6640), .S(n4070), .Z(n6653) );
  CMX2X1 U15429 ( .A0(n6641), .A1(n6653), .S(n3771), .Z(n6666) );
  CMXI2X1 U15430 ( .A0(n6642), .A1(n6666), .S(n3487), .Z(N2194) );
  CMX2X1 U15431 ( .A0(mem_data1[133]), .A1(mem_data1[134]), .S(n3862), .Z(
        n6649) );
  CMXI2X1 U15432 ( .A0(n6649), .A1(n6643), .S(n4070), .Z(n6656) );
  CMX2X1 U15433 ( .A0(n6644), .A1(n6656), .S(n3772), .Z(n6669) );
  CMXI2X1 U15434 ( .A0(n6645), .A1(n6669), .S(n3487), .Z(N2195) );
  CMX2X1 U15435 ( .A0(mem_data1[13]), .A1(mem_data1[14]), .S(n3878), .Z(n6712)
         );
  CMX2X1 U15436 ( .A0(mem_data1[11]), .A1(mem_data1[12]), .S(n3877), .Z(n6923)
         );
  CMXI2X1 U15437 ( .A0(n6712), .A1(n6923), .S(n4070), .Z(n8932) );
  CMX2X1 U15438 ( .A0(mem_data1[17]), .A1(mem_data1[18]), .S(n3863), .Z(n6714)
         );
  CMX2X1 U15439 ( .A0(mem_data1[15]), .A1(mem_data1[16]), .S(n3880), .Z(n6713)
         );
  CMXI2X1 U15440 ( .A0(n6714), .A1(n6713), .S(n4070), .Z(n6784) );
  CMX2X1 U15441 ( .A0(n8932), .A1(n6784), .S(n3773), .Z(n7598) );
  CMX2X1 U15442 ( .A0(mem_data1[21]), .A1(mem_data1[22]), .S(n3881), .Z(n6716)
         );
  CMX2X1 U15443 ( .A0(mem_data1[19]), .A1(mem_data1[20]), .S(n3862), .Z(n6715)
         );
  CMXI2X1 U15444 ( .A0(n6716), .A1(n6715), .S(n4070), .Z(n6783) );
  CMX2X1 U15445 ( .A0(mem_data1[25]), .A1(mem_data1[26]), .S(n3863), .Z(n6718)
         );
  CMX2X1 U15446 ( .A0(mem_data1[23]), .A1(mem_data1[24]), .S(n3871), .Z(n6717)
         );
  CMXI2X1 U15447 ( .A0(n6718), .A1(n6717), .S(n4070), .Z(n6786) );
  CMX2X1 U15448 ( .A0(n6783), .A1(n6786), .S(n3774), .Z(n6920) );
  CMXI2X1 U15449 ( .A0(n7598), .A1(n6920), .S(n3487), .Z(N2087) );
  CMX2X1 U15450 ( .A0(mem_data1[134]), .A1(mem_data1[135]), .S(n3862), .Z(
        n6652) );
  CMXI2X1 U15451 ( .A0(n6652), .A1(n6646), .S(n4070), .Z(n6659) );
  CMX2X1 U15452 ( .A0(n6647), .A1(n6659), .S(n3775), .Z(n6672) );
  CMXI2X1 U15453 ( .A0(n6648), .A1(n6672), .S(n3487), .Z(N2196) );
  CMX2X1 U15454 ( .A0(mem_data1[135]), .A1(mem_data1[136]), .S(n3863), .Z(
        n6655) );
  CMXI2X1 U15455 ( .A0(n6655), .A1(n6649), .S(n4070), .Z(n6662) );
  CMX2X1 U15456 ( .A0(n6650), .A1(n6662), .S(n3776), .Z(n6675) );
  CMXI2X1 U15457 ( .A0(n6651), .A1(n6675), .S(n3487), .Z(N2197) );
  CMX2X1 U15458 ( .A0(mem_data1[136]), .A1(mem_data1[137]), .S(n3878), .Z(
        n6658) );
  CMXI2X1 U15459 ( .A0(n6658), .A1(n6652), .S(n4070), .Z(n6665) );
  CMX2X1 U15460 ( .A0(n6653), .A1(n6665), .S(n3777), .Z(n6684) );
  CMXI2X1 U15461 ( .A0(n6654), .A1(n6684), .S(n3487), .Z(N2198) );
  CMX2X1 U15462 ( .A0(mem_data1[137]), .A1(mem_data1[138]), .S(n3879), .Z(
        n6661) );
  CMXI2X1 U15463 ( .A0(n6661), .A1(n6655), .S(n4070), .Z(n6668) );
  CMX2X1 U15464 ( .A0(n6656), .A1(n6668), .S(n3790), .Z(n6687) );
  CMXI2X1 U15465 ( .A0(n6657), .A1(n6687), .S(n3487), .Z(N2199) );
  CMX2X1 U15466 ( .A0(mem_data1[138]), .A1(mem_data1[139]), .S(n3864), .Z(
        n6664) );
  CMXI2X1 U15467 ( .A0(n6664), .A1(n6658), .S(n4069), .Z(n6671) );
  CMX2X1 U15468 ( .A0(n6659), .A1(n6671), .S(n3791), .Z(n6690) );
  CMXI2X1 U15469 ( .A0(n6660), .A1(n6690), .S(n3487), .Z(N2200) );
  CMX2X1 U15470 ( .A0(mem_data1[139]), .A1(mem_data1[140]), .S(n3865), .Z(
        n6667) );
  CMXI2X1 U15471 ( .A0(n6667), .A1(n6661), .S(n4069), .Z(n6674) );
  CMX2X1 U15472 ( .A0(n6662), .A1(n6674), .S(n4367), .Z(n6693) );
  CMXI2X1 U15473 ( .A0(n6663), .A1(n6693), .S(n3486), .Z(N2201) );
  CMX2X1 U15474 ( .A0(mem_data1[140]), .A1(mem_data1[141]), .S(n3866), .Z(
        n6670) );
  CMXI2X1 U15475 ( .A0(n6670), .A1(n6664), .S(n4069), .Z(n6683) );
  CMX2X1 U15476 ( .A0(n6665), .A1(n6683), .S(n3790), .Z(n6696) );
  CMXI2X1 U15477 ( .A0(n6666), .A1(n6696), .S(n3486), .Z(N2202) );
  CMX2X1 U15478 ( .A0(mem_data1[141]), .A1(mem_data1[142]), .S(n3867), .Z(
        n6673) );
  CMXI2X1 U15479 ( .A0(n6673), .A1(n6667), .S(n4069), .Z(n6686) );
  CMX2X1 U15480 ( .A0(n6668), .A1(n6686), .S(n3793), .Z(n6699) );
  CMXI2X1 U15481 ( .A0(n6669), .A1(n6699), .S(n3486), .Z(N2203) );
  CMX2X1 U15482 ( .A0(mem_data1[142]), .A1(mem_data1[143]), .S(n3877), .Z(
        n6682) );
  CMXI2X1 U15483 ( .A0(n6682), .A1(n6670), .S(n4069), .Z(n6689) );
  CMX2X1 U15484 ( .A0(n6671), .A1(n6689), .S(n3794), .Z(n6702) );
  CMXI2X1 U15485 ( .A0(n6672), .A1(n6702), .S(n3486), .Z(N2204) );
  CMX2X1 U15486 ( .A0(mem_data1[143]), .A1(mem_data1[144]), .S(n3878), .Z(
        n6685) );
  CMXI2X1 U15487 ( .A0(n6685), .A1(n6673), .S(n4069), .Z(n6692) );
  CMX2X1 U15488 ( .A0(n6674), .A1(n6692), .S(n3795), .Z(n6705) );
  CMXI2X1 U15489 ( .A0(n6675), .A1(n6705), .S(n3486), .Z(N2205) );
  CMXI2X1 U15490 ( .A0(n6677), .A1(n6676), .S(n4069), .Z(n6818) );
  CMX2X1 U15491 ( .A0(n6678), .A1(n6818), .S(n3796), .Z(n7932) );
  CMXI2X1 U15492 ( .A0(n6680), .A1(n6679), .S(n4069), .Z(n6817) );
  CMX2X1 U15493 ( .A0(mem_data1[26]), .A1(mem_data1[27]), .S(n3879), .Z(n6751)
         );
  CMXI2X1 U15494 ( .A0(n6751), .A1(n6681), .S(n4069), .Z(n6820) );
  CMX2X1 U15495 ( .A0(n6817), .A1(n6820), .S(n3797), .Z(n6958) );
  CMXI2X1 U15496 ( .A0(n7932), .A1(n6958), .S(n3486), .Z(N2088) );
  CMX2X1 U15497 ( .A0(mem_data1[144]), .A1(mem_data1[145]), .S(n3880), .Z(
        n6688) );
  CMXI2X1 U15498 ( .A0(n6688), .A1(n6682), .S(n4069), .Z(n6695) );
  CMX2X1 U15499 ( .A0(n6683), .A1(n6695), .S(n4364), .Z(n6708) );
  CMXI2X1 U15500 ( .A0(n6684), .A1(n6708), .S(n3486), .Z(N2206) );
  CMX2X1 U15501 ( .A0(mem_data1[145]), .A1(mem_data1[146]), .S(n3872), .Z(
        n6691) );
  CMXI2X1 U15502 ( .A0(n6691), .A1(n6685), .S(n4069), .Z(n6698) );
  CMX2X1 U15503 ( .A0(n6686), .A1(n6698), .S(n4364), .Z(n6711) );
  CMXI2X1 U15504 ( .A0(n6687), .A1(n6711), .S(n3486), .Z(N2207) );
  CMX2X1 U15505 ( .A0(mem_data1[146]), .A1(mem_data1[147]), .S(n3880), .Z(
        n6694) );
  CMXI2X1 U15506 ( .A0(n6694), .A1(n6688), .S(n4069), .Z(n6701) );
  CMX2X1 U15507 ( .A0(n6689), .A1(n6701), .S(n4364), .Z(n6721) );
  CMXI2X1 U15508 ( .A0(n6690), .A1(n6721), .S(n3486), .Z(N2208) );
  CMX2X1 U15509 ( .A0(mem_data1[147]), .A1(mem_data1[148]), .S(n3881), .Z(
        n6697) );
  CMXI2X1 U15510 ( .A0(n6697), .A1(n6691), .S(n4069), .Z(n6704) );
  CMX2X1 U15511 ( .A0(n6692), .A1(n6704), .S(n4364), .Z(n6724) );
  CMXI2X1 U15512 ( .A0(n6693), .A1(n6724), .S(n3486), .Z(N2209) );
  CMX2X1 U15513 ( .A0(mem_data1[148]), .A1(mem_data1[149]), .S(n3862), .Z(
        n6700) );
  CMXI2X1 U15514 ( .A0(n6700), .A1(n6694), .S(n4069), .Z(n6707) );
  CMX2X1 U15515 ( .A0(n6695), .A1(n6707), .S(n4364), .Z(n6727) );
  CMXI2X1 U15516 ( .A0(n6696), .A1(n6727), .S(n3489), .Z(N2210) );
  CMX2X1 U15517 ( .A0(mem_data1[149]), .A1(mem_data1[150]), .S(n3863), .Z(
        n6703) );
  CMXI2X1 U15518 ( .A0(n6703), .A1(n6697), .S(n4069), .Z(n6710) );
  CMX2X1 U15519 ( .A0(n6698), .A1(n6710), .S(n4364), .Z(n6730) );
  CMXI2X1 U15520 ( .A0(n6699), .A1(n6730), .S(n3489), .Z(N2211) );
  CMX2X1 U15521 ( .A0(mem_data1[150]), .A1(mem_data1[151]), .S(n3864), .Z(
        n6706) );
  CMXI2X1 U15522 ( .A0(n6706), .A1(n6700), .S(n4069), .Z(n6720) );
  CMX2X1 U15523 ( .A0(n6701), .A1(n6720), .S(n4364), .Z(n6733) );
  CMXI2X1 U15524 ( .A0(n6702), .A1(n6733), .S(n3489), .Z(N2212) );
  CMX2X1 U15525 ( .A0(mem_data1[151]), .A1(mem_data1[152]), .S(n3865), .Z(
        n6709) );
  CMXI2X1 U15526 ( .A0(n6709), .A1(n6703), .S(n4068), .Z(n6723) );
  CMX2X1 U15527 ( .A0(n6704), .A1(n6723), .S(n4364), .Z(n6736) );
  CMXI2X1 U15528 ( .A0(n6705), .A1(n6736), .S(n3489), .Z(N2213) );
  CMX2X1 U15529 ( .A0(mem_data1[152]), .A1(mem_data1[153]), .S(n3866), .Z(
        n6719) );
  CMXI2X1 U15530 ( .A0(n6719), .A1(n6706), .S(n4068), .Z(n6726) );
  CMX2X1 U15531 ( .A0(n6707), .A1(n6726), .S(n4364), .Z(n6739) );
  CMXI2X1 U15532 ( .A0(n6708), .A1(n6739), .S(n3488), .Z(N2214) );
  CMX2X1 U15533 ( .A0(mem_data1[153]), .A1(mem_data1[154]), .S(n3864), .Z(
        n6722) );
  CMXI2X1 U15534 ( .A0(n6722), .A1(n6709), .S(n4068), .Z(n6729) );
  CMX2X1 U15535 ( .A0(n6710), .A1(n6729), .S(n4364), .Z(n6742) );
  CMXI2X1 U15536 ( .A0(n6711), .A1(n6742), .S(n3488), .Z(N2215) );
  CMXI2X1 U15537 ( .A0(n6713), .A1(n6712), .S(n4068), .Z(n6924) );
  CMXI2X1 U15538 ( .A0(n6715), .A1(n6714), .S(n4068), .Z(n6852) );
  CMX2X1 U15539 ( .A0(n6924), .A1(n6852), .S(n4364), .Z(n8266) );
  CMXI2X1 U15540 ( .A0(n6717), .A1(n6716), .S(n4068), .Z(n6851) );
  CMX2X1 U15541 ( .A0(mem_data1[27]), .A1(mem_data1[28]), .S(n3865), .Z(n6785)
         );
  CMXI2X1 U15542 ( .A0(n6785), .A1(n6718), .S(n4068), .Z(n6854) );
  CMX2X1 U15543 ( .A0(n6851), .A1(n6854), .S(n4363), .Z(n6991) );
  CMXI2X1 U15544 ( .A0(n8266), .A1(n6991), .S(n3488), .Z(N2089) );
  CMX2X1 U15545 ( .A0(mem_data1[154]), .A1(mem_data1[155]), .S(n3868), .Z(
        n6725) );
  CMXI2X1 U15546 ( .A0(n6725), .A1(n6719), .S(n4068), .Z(n6732) );
  CMX2X1 U15547 ( .A0(n6720), .A1(n6732), .S(n4363), .Z(n6745) );
  CMXI2X1 U15548 ( .A0(n6721), .A1(n6745), .S(n3488), .Z(N2216) );
  CMX2X1 U15549 ( .A0(mem_data1[155]), .A1(mem_data1[156]), .S(n3868), .Z(
        n6728) );
  CMXI2X1 U15550 ( .A0(n6728), .A1(n6722), .S(n4068), .Z(n6735) );
  CMX2X1 U15551 ( .A0(n6723), .A1(n6735), .S(n4363), .Z(n6748) );
  CMXI2X1 U15552 ( .A0(n6724), .A1(n6748), .S(n3488), .Z(N2217) );
  CMX2X1 U15553 ( .A0(mem_data1[156]), .A1(mem_data1[157]), .S(n3869), .Z(
        n6731) );
  CMXI2X1 U15554 ( .A0(n6731), .A1(n6725), .S(n4068), .Z(n6738) );
  CMX2X1 U15555 ( .A0(n6726), .A1(n6738), .S(n4363), .Z(n6755) );
  CMXI2X1 U15556 ( .A0(n6727), .A1(n6755), .S(n3488), .Z(N2218) );
  CMX2X1 U15557 ( .A0(mem_data1[157]), .A1(mem_data1[158]), .S(n3870), .Z(
        n6734) );
  CMXI2X1 U15558 ( .A0(n6734), .A1(n6728), .S(n4068), .Z(n6741) );
  CMX2X1 U15559 ( .A0(n6729), .A1(n6741), .S(n4363), .Z(n6758) );
  CMXI2X1 U15560 ( .A0(n6730), .A1(n6758), .S(n3488), .Z(N2219) );
  CMX2X1 U15561 ( .A0(mem_data1[158]), .A1(mem_data1[159]), .S(n3871), .Z(
        n6737) );
  CMXI2X1 U15562 ( .A0(n6737), .A1(n6731), .S(n4068), .Z(n6744) );
  CMX2X1 U15563 ( .A0(n6732), .A1(n6744), .S(n4363), .Z(n6761) );
  CMXI2X1 U15564 ( .A0(n6733), .A1(n6761), .S(n3488), .Z(N2220) );
  CMX2X1 U15565 ( .A0(mem_data1[159]), .A1(mem_data1[160]), .S(n3881), .Z(
        n6740) );
  CMXI2X1 U15566 ( .A0(n6740), .A1(n6734), .S(n4068), .Z(n6747) );
  CMX2X1 U15567 ( .A0(n6735), .A1(n6747), .S(n4363), .Z(n6764) );
  CMXI2X1 U15568 ( .A0(n6736), .A1(n6764), .S(n3488), .Z(N2221) );
  CMX2X1 U15569 ( .A0(mem_data1[160]), .A1(mem_data1[161]), .S(n3862), .Z(
        n6743) );
  CMXI2X1 U15570 ( .A0(n6743), .A1(n6737), .S(n4068), .Z(n6754) );
  CMX2X1 U15571 ( .A0(n6738), .A1(n6754), .S(n4363), .Z(n6767) );
  CMXI2X1 U15572 ( .A0(n6739), .A1(n6767), .S(n3488), .Z(N2222) );
  CMX2X1 U15573 ( .A0(mem_data1[161]), .A1(mem_data1[162]), .S(n3863), .Z(
        n6746) );
  CMXI2X1 U15574 ( .A0(n6746), .A1(n6740), .S(n4068), .Z(n6757) );
  CMX2X1 U15575 ( .A0(n6741), .A1(n6757), .S(n4363), .Z(n6770) );
  CMXI2X1 U15576 ( .A0(n6742), .A1(n6770), .S(n3488), .Z(N2223) );
  CMX2X1 U15577 ( .A0(mem_data1[162]), .A1(mem_data1[163]), .S(n3864), .Z(
        n6753) );
  CMXI2X1 U15578 ( .A0(n6753), .A1(n6743), .S(n4068), .Z(n6760) );
  CMX2X1 U15579 ( .A0(n6744), .A1(n6760), .S(n4363), .Z(n6773) );
  CMXI2X1 U15580 ( .A0(n6745), .A1(n6773), .S(n3487), .Z(N2224) );
  CMX2X1 U15581 ( .A0(mem_data1[163]), .A1(mem_data1[164]), .S(n3873), .Z(
        n6756) );
  CMXI2X1 U15582 ( .A0(n6756), .A1(n6746), .S(n4067), .Z(n6763) );
  CMX2X1 U15583 ( .A0(n6747), .A1(n6763), .S(n4363), .Z(n6776) );
  CMXI2X1 U15584 ( .A0(n6748), .A1(n6776), .S(n3487), .Z(N2225) );
  CMX2X1 U15585 ( .A0(n6750), .A1(n6749), .S(n4362), .Z(n8600) );
  CMX2X1 U15586 ( .A0(mem_data1[28]), .A1(mem_data1[29]), .S(n3869), .Z(n6819)
         );
  CMXI2X1 U15587 ( .A0(n6819), .A1(n6751), .S(n4067), .Z(n6886) );
  CMX2X1 U15588 ( .A0(n6752), .A1(n6886), .S(n4362), .Z(n7024) );
  CMXI2X1 U15589 ( .A0(n8600), .A1(n7024), .S(n3487), .Z(N2090) );
  CMX2X1 U15590 ( .A0(mem_data1[164]), .A1(mem_data1[165]), .S(n3870), .Z(
        n6759) );
  CMXI2X1 U15591 ( .A0(n6759), .A1(n6753), .S(n4067), .Z(n6766) );
  CMX2X1 U15592 ( .A0(n6754), .A1(n6766), .S(n4362), .Z(n6779) );
  CMXI2X1 U15593 ( .A0(n6755), .A1(n6779), .S(n3491), .Z(N2226) );
  CMX2X1 U15594 ( .A0(mem_data1[165]), .A1(mem_data1[166]), .S(n3871), .Z(
        n6762) );
  CMXI2X1 U15595 ( .A0(n6762), .A1(n6756), .S(n4067), .Z(n6769) );
  CMX2X1 U15596 ( .A0(n6757), .A1(n6769), .S(n4362), .Z(n6782) );
  CMXI2X1 U15597 ( .A0(n6758), .A1(n6782), .S(n3490), .Z(N2227) );
  CMX2X1 U15598 ( .A0(mem_data1[166]), .A1(mem_data1[167]), .S(n3872), .Z(
        n6765) );
  CMXI2X1 U15599 ( .A0(n6765), .A1(n6759), .S(n4067), .Z(n6772) );
  CMX2X1 U15600 ( .A0(n6760), .A1(n6772), .S(n4362), .Z(n6789) );
  CMXI2X1 U15601 ( .A0(n6761), .A1(n6789), .S(n3490), .Z(N2228) );
  CMX2X1 U15602 ( .A0(mem_data1[167]), .A1(mem_data1[168]), .S(n3873), .Z(
        n6768) );
  CMXI2X1 U15603 ( .A0(n6768), .A1(n6762), .S(n4067), .Z(n6775) );
  CMX2X1 U15604 ( .A0(n6763), .A1(n6775), .S(n4362), .Z(n6792) );
  CMXI2X1 U15605 ( .A0(n6764), .A1(n6792), .S(n3490), .Z(N2229) );
  CMX2X1 U15606 ( .A0(mem_data1[168]), .A1(mem_data1[169]), .S(n3874), .Z(
        n6771) );
  CMXI2X1 U15607 ( .A0(n6771), .A1(n6765), .S(n4067), .Z(n6778) );
  CMX2X1 U15608 ( .A0(n6766), .A1(n6778), .S(n4362), .Z(n6795) );
  CMXI2X1 U15609 ( .A0(n6767), .A1(n6795), .S(n3490), .Z(N2230) );
  CMX2X1 U15610 ( .A0(mem_data1[169]), .A1(mem_data1[170]), .S(n3875), .Z(
        n6774) );
  CMXI2X1 U15611 ( .A0(n6774), .A1(n6768), .S(n4067), .Z(n6781) );
  CMX2X1 U15612 ( .A0(n6769), .A1(n6781), .S(n4362), .Z(n6798) );
  CMXI2X1 U15613 ( .A0(n6770), .A1(n6798), .S(n3490), .Z(N2231) );
  CMX2X1 U15614 ( .A0(mem_data1[170]), .A1(mem_data1[171]), .S(n3866), .Z(
        n6777) );
  CMXI2X1 U15615 ( .A0(n6777), .A1(n6771), .S(n4067), .Z(n6788) );
  CMX2X1 U15616 ( .A0(n6772), .A1(n6788), .S(n4362), .Z(n6801) );
  CMXI2X1 U15617 ( .A0(n6773), .A1(n6801), .S(n3490), .Z(N2232) );
  CMX2X1 U15618 ( .A0(mem_data1[171]), .A1(mem_data1[172]), .S(n3867), .Z(
        n6780) );
  CMXI2X1 U15619 ( .A0(n6780), .A1(n6774), .S(n4067), .Z(n6791) );
  CMX2X1 U15620 ( .A0(n6775), .A1(n6791), .S(n4362), .Z(n6804) );
  CMXI2X1 U15621 ( .A0(n6776), .A1(n6804), .S(n3490), .Z(N2233) );
  CMX2X1 U15622 ( .A0(mem_data1[172]), .A1(mem_data1[173]), .S(n3876), .Z(
        n6787) );
  CMXI2X1 U15623 ( .A0(n6787), .A1(n6777), .S(n4067), .Z(n6794) );
  CMX2X1 U15624 ( .A0(n6778), .A1(n6794), .S(n4361), .Z(n6807) );
  CMXI2X1 U15625 ( .A0(n6779), .A1(n6807), .S(n3490), .Z(N2234) );
  CMX2X1 U15626 ( .A0(mem_data1[173]), .A1(mem_data1[174]), .S(n3877), .Z(
        n6790) );
  CMXI2X1 U15627 ( .A0(n6790), .A1(n6780), .S(n4067), .Z(n6797) );
  CMX2X1 U15628 ( .A0(n6781), .A1(n6797), .S(n4361), .Z(n6810) );
  CMXI2X1 U15629 ( .A0(n6782), .A1(n6810), .S(n3490), .Z(N2235) );
  CMX2X1 U15630 ( .A0(n6784), .A1(n6783), .S(n4361), .Z(n8934) );
  CMX2X1 U15631 ( .A0(mem_data1[29]), .A1(mem_data1[30]), .S(n3872), .Z(n6853)
         );
  CMXI2X1 U15632 ( .A0(n6853), .A1(n6785), .S(n4067), .Z(n6919) );
  CMX2X1 U15633 ( .A0(n6786), .A1(n6919), .S(n4361), .Z(n7057) );
  CMXI2X1 U15634 ( .A0(n8934), .A1(n7057), .S(n3490), .Z(N2091) );
  CMX2X1 U15635 ( .A0(mem_data1[174]), .A1(mem_data1[175]), .S(n3873), .Z(
        n6793) );
  CMXI2X1 U15636 ( .A0(n6793), .A1(n6787), .S(n4067), .Z(n6800) );
  CMX2X1 U15637 ( .A0(n6788), .A1(n6800), .S(n4361), .Z(n6813) );
  CMXI2X1 U15638 ( .A0(n6789), .A1(n6813), .S(n3490), .Z(N2236) );
  CMX2X1 U15639 ( .A0(mem_data1[175]), .A1(mem_data1[176]), .S(n3874), .Z(
        n6796) );
  CMXI2X1 U15640 ( .A0(n6796), .A1(n6790), .S(n4067), .Z(n6803) );
  CMX2X1 U15641 ( .A0(n6791), .A1(n6803), .S(n4361), .Z(n6816) );
  CMXI2X1 U15642 ( .A0(n6792), .A1(n6816), .S(n3489), .Z(N2237) );
  CMX2X1 U15643 ( .A0(mem_data1[176]), .A1(mem_data1[177]), .S(n3875), .Z(
        n6799) );
  CMXI2X1 U15644 ( .A0(n6799), .A1(n6793), .S(n4067), .Z(n6806) );
  CMX2X1 U15645 ( .A0(n6794), .A1(n6806), .S(n4361), .Z(n6823) );
  CMXI2X1 U15646 ( .A0(n6795), .A1(n6823), .S(n3489), .Z(N2238) );
  CMX2X1 U15647 ( .A0(mem_data1[177]), .A1(mem_data1[178]), .S(n3865), .Z(
        n6802) );
  CMXI2X1 U15648 ( .A0(n6802), .A1(n6796), .S(n4066), .Z(n6809) );
  CMX2X1 U15649 ( .A0(n6797), .A1(n6809), .S(n4361), .Z(n6826) );
  CMXI2X1 U15650 ( .A0(n6798), .A1(n6826), .S(n3489), .Z(N2239) );
  CMX2X1 U15651 ( .A0(mem_data1[178]), .A1(mem_data1[179]), .S(n3866), .Z(
        n6805) );
  CMXI2X1 U15652 ( .A0(n6805), .A1(n6799), .S(n4066), .Z(n6812) );
  CMX2X1 U15653 ( .A0(n6800), .A1(n6812), .S(n4361), .Z(n6829) );
  CMXI2X1 U15654 ( .A0(n6801), .A1(n6829), .S(n3489), .Z(N2240) );
  CMX2X1 U15655 ( .A0(mem_data1[179]), .A1(mem_data1[180]), .S(n3867), .Z(
        n6808) );
  CMXI2X1 U15656 ( .A0(n6808), .A1(n6802), .S(n4066), .Z(n6815) );
  CMX2X1 U15657 ( .A0(n6803), .A1(n6815), .S(n4361), .Z(n6832) );
  CMXI2X1 U15658 ( .A0(n6804), .A1(n6832), .S(n3489), .Z(N2241) );
  CMX2X1 U15659 ( .A0(mem_data1[180]), .A1(mem_data1[181]), .S(n3868), .Z(
        n6811) );
  CMXI2X1 U15660 ( .A0(n6811), .A1(n6805), .S(n4066), .Z(n6822) );
  CMX2X1 U15661 ( .A0(n6806), .A1(n6822), .S(n4361), .Z(n6835) );
  CMXI2X1 U15662 ( .A0(n6807), .A1(n6835), .S(n3489), .Z(N2242) );
  CMX2X1 U15663 ( .A0(mem_data1[181]), .A1(mem_data1[182]), .S(n3874), .Z(
        n6814) );
  CMXI2X1 U15664 ( .A0(n6814), .A1(n6808), .S(n4066), .Z(n6825) );
  CMX2X1 U15665 ( .A0(n6809), .A1(n6825), .S(n4360), .Z(n6838) );
  CMXI2X1 U15666 ( .A0(n6810), .A1(n6838), .S(n3492), .Z(N2243) );
  CMX2X1 U15667 ( .A0(mem_data1[182]), .A1(mem_data1[183]), .S(n3878), .Z(
        n6821) );
  CMXI2X1 U15668 ( .A0(n6821), .A1(n6811), .S(n4066), .Z(n6828) );
  CMX2X1 U15669 ( .A0(n6812), .A1(n6828), .S(n4360), .Z(n6841) );
  CMXI2X1 U15670 ( .A0(n6813), .A1(n6841), .S(n3492), .Z(N2244) );
  CMX2X1 U15671 ( .A0(mem_data1[183]), .A1(mem_data1[184]), .S(n3879), .Z(
        n6824) );
  CMXI2X1 U15672 ( .A0(n6824), .A1(n6814), .S(n4066), .Z(n6831) );
  CMX2X1 U15673 ( .A0(n6815), .A1(n6831), .S(n4360), .Z(n6844) );
  CMXI2X1 U15674 ( .A0(n6816), .A1(n6844), .S(n3492), .Z(N2245) );
  CMX2X1 U15675 ( .A0(n6818), .A1(n6817), .S(n4360), .Z(n9268) );
  CMX2X1 U15676 ( .A0(mem_data1[30]), .A1(mem_data1[31]), .S(n3880), .Z(n6885)
         );
  CMXI2X1 U15677 ( .A0(n6885), .A1(n6819), .S(n4066), .Z(n6957) );
  CMX2X1 U15678 ( .A0(n6820), .A1(n6957), .S(n4360), .Z(n7090) );
  CMXI2X1 U15679 ( .A0(n9268), .A1(n7090), .S(n3492), .Z(N2092) );
  CMX2X1 U15680 ( .A0(mem_data1[184]), .A1(mem_data1[185]), .S(n3881), .Z(
        n6827) );
  CMXI2X1 U15681 ( .A0(n6827), .A1(n6821), .S(n4066), .Z(n6834) );
  CMX2X1 U15682 ( .A0(n6822), .A1(n6834), .S(n4360), .Z(n6847) );
  CMXI2X1 U15683 ( .A0(n6823), .A1(n6847), .S(n3492), .Z(N2246) );
  CMX2X1 U15684 ( .A0(mem_data1[185]), .A1(mem_data1[186]), .S(n3862), .Z(
        n6830) );
  CMXI2X1 U15685 ( .A0(n6830), .A1(n6824), .S(n4066), .Z(n6837) );
  CMX2X1 U15686 ( .A0(n6825), .A1(n6837), .S(n4360), .Z(n6850) );
  CMXI2X1 U15687 ( .A0(n6826), .A1(n6850), .S(n3492), .Z(N2247) );
  CMX2X1 U15688 ( .A0(mem_data1[186]), .A1(mem_data1[187]), .S(n3863), .Z(
        n6833) );
  CMXI2X1 U15689 ( .A0(n6833), .A1(n6827), .S(n4066), .Z(n6840) );
  CMX2X1 U15690 ( .A0(n6828), .A1(n6840), .S(n4360), .Z(n6857) );
  CMXI2X1 U15691 ( .A0(n6829), .A1(n6857), .S(n3492), .Z(N2248) );
  CMX2X1 U15692 ( .A0(mem_data1[187]), .A1(mem_data1[188]), .S(n3864), .Z(
        n6836) );
  CMXI2X1 U15693 ( .A0(n6836), .A1(n6830), .S(n4066), .Z(n6843) );
  CMX2X1 U15694 ( .A0(n6831), .A1(n6843), .S(n4360), .Z(n6860) );
  CMXI2X1 U15695 ( .A0(n6832), .A1(n6860), .S(n3491), .Z(N2249) );
  CMX2X1 U15696 ( .A0(mem_data1[188]), .A1(mem_data1[189]), .S(n3868), .Z(
        n6839) );
  CMXI2X1 U15697 ( .A0(n6839), .A1(n6833), .S(n4066), .Z(n6846) );
  CMX2X1 U15698 ( .A0(n6834), .A1(n6846), .S(n4360), .Z(n6863) );
  CMXI2X1 U15699 ( .A0(n6835), .A1(n6863), .S(n3491), .Z(N2250) );
  CMX2X1 U15700 ( .A0(mem_data1[189]), .A1(mem_data1[190]), .S(n3869), .Z(
        n6842) );
  CMXI2X1 U15701 ( .A0(n6842), .A1(n6836), .S(n4066), .Z(n6849) );
  CMX2X1 U15702 ( .A0(n6837), .A1(n6849), .S(n4360), .Z(n6866) );
  CMXI2X1 U15703 ( .A0(n6838), .A1(n6866), .S(n3491), .Z(N2251) );
  CMX2X1 U15704 ( .A0(mem_data1[190]), .A1(mem_data1[191]), .S(n3865), .Z(
        n6845) );
  CMXI2X1 U15705 ( .A0(n6845), .A1(n6839), .S(n4066), .Z(n6856) );
  CMX2X1 U15706 ( .A0(n6840), .A1(n6856), .S(n4359), .Z(n6869) );
  CMXI2X1 U15707 ( .A0(n6841), .A1(n6869), .S(n3491), .Z(N2252) );
  CMX2X1 U15708 ( .A0(mem_data1[191]), .A1(mem_data1[192]), .S(n3866), .Z(
        n6848) );
  CMXI2X1 U15709 ( .A0(n6848), .A1(n6842), .S(n4066), .Z(n6859) );
  CMX2X1 U15710 ( .A0(n6843), .A1(n6859), .S(n4359), .Z(n6872) );
  CMXI2X1 U15711 ( .A0(n6844), .A1(n6872), .S(n3491), .Z(N2253) );
  CMX2X1 U15712 ( .A0(mem_data1[192]), .A1(mem_data1[193]), .S(n3876), .Z(
        n6855) );
  CMXI2X1 U15713 ( .A0(n6855), .A1(n6845), .S(n4065), .Z(n6862) );
  CMX2X1 U15714 ( .A0(n6846), .A1(n6862), .S(n4359), .Z(n6875) );
  CMXI2X1 U15715 ( .A0(n6847), .A1(n6875), .S(n3491), .Z(N2254) );
  CMX2X1 U15716 ( .A0(mem_data1[193]), .A1(mem_data1[194]), .S(n3877), .Z(
        n6858) );
  CMXI2X1 U15717 ( .A0(n6858), .A1(n6848), .S(n4065), .Z(n6865) );
  CMX2X1 U15718 ( .A0(n6849), .A1(n6865), .S(n4359), .Z(n6878) );
  CMXI2X1 U15719 ( .A0(n6850), .A1(n6878), .S(n3491), .Z(N2255) );
  CMX2X1 U15720 ( .A0(n6852), .A1(n6851), .S(n4359), .Z(n9586) );
  CMX2X1 U15721 ( .A0(mem_data1[31]), .A1(mem_data1[32]), .S(n3878), .Z(n6918)
         );
  CMXI2X1 U15722 ( .A0(n6918), .A1(n6853), .S(n4065), .Z(n6990) );
  CMX2X1 U15723 ( .A0(n6854), .A1(n6990), .S(n4359), .Z(n7123) );
  CMXI2X1 U15724 ( .A0(n9586), .A1(n7123), .S(n3491), .Z(N2093) );
  CMX2X1 U15725 ( .A0(mem_data1[194]), .A1(mem_data1[195]), .S(n3879), .Z(
        n6861) );
  CMXI2X1 U15726 ( .A0(n6861), .A1(n6855), .S(n4065), .Z(n6868) );
  CMX2X1 U15727 ( .A0(n6856), .A1(n6868), .S(n4359), .Z(n6881) );
  CMXI2X1 U15728 ( .A0(n6857), .A1(n6881), .S(n3491), .Z(N2256) );
  CMX2X1 U15729 ( .A0(mem_data1[195]), .A1(mem_data1[196]), .S(n3869), .Z(
        n6864) );
  CMXI2X1 U15730 ( .A0(n6864), .A1(n6858), .S(n4065), .Z(n6871) );
  CMX2X1 U15731 ( .A0(n6859), .A1(n6871), .S(n4359), .Z(n6884) );
  CMXI2X1 U15732 ( .A0(n6860), .A1(n6884), .S(n3491), .Z(N2257) );
  CMX2X1 U15733 ( .A0(mem_data1[196]), .A1(mem_data1[197]), .S(n3870), .Z(
        n6867) );
  CMXI2X1 U15734 ( .A0(n6867), .A1(n6861), .S(n4065), .Z(n6874) );
  CMX2X1 U15735 ( .A0(n6862), .A1(n6874), .S(n4359), .Z(n6890) );
  CMXI2X1 U15736 ( .A0(n6863), .A1(n6890), .S(n3494), .Z(N2258) );
  CMX2X1 U15737 ( .A0(mem_data1[197]), .A1(mem_data1[198]), .S(n3871), .Z(
        n6870) );
  CMXI2X1 U15738 ( .A0(n6870), .A1(n6864), .S(n4065), .Z(n6877) );
  CMX2X1 U15739 ( .A0(n6865), .A1(n6877), .S(n4359), .Z(n6893) );
  CMXI2X1 U15740 ( .A0(n6866), .A1(n6893), .S(n3494), .Z(N2259) );
  CMX2X1 U15741 ( .A0(mem_data1[198]), .A1(mem_data1[199]), .S(n3872), .Z(
        n6873) );
  CMXI2X1 U15742 ( .A0(n6873), .A1(n6867), .S(n4065), .Z(n6880) );
  CMX2X1 U15743 ( .A0(n6868), .A1(n6880), .S(n4359), .Z(n6896) );
  CMXI2X1 U15744 ( .A0(n6869), .A1(n6896), .S(n3494), .Z(N2260) );
  CMX2X1 U15745 ( .A0(mem_data1[199]), .A1(mem_data1[200]), .S(n3875), .Z(
        n6876) );
  CMXI2X1 U15746 ( .A0(n6876), .A1(n6870), .S(n4065), .Z(n6883) );
  CMX2X1 U15747 ( .A0(n6871), .A1(n6883), .S(n4358), .Z(n6899) );
  CMXI2X1 U15748 ( .A0(n6872), .A1(n6899), .S(n3494), .Z(N2261) );
  CMX2X1 U15749 ( .A0(mem_data1[200]), .A1(mem_data1[201]), .S(n3867), .Z(
        n6879) );
  CMXI2X1 U15750 ( .A0(n6879), .A1(n6873), .S(n4065), .Z(n6889) );
  CMX2X1 U15751 ( .A0(n6874), .A1(n6889), .S(n4358), .Z(n6902) );
  CMXI2X1 U15752 ( .A0(n6875), .A1(n6902), .S(n3493), .Z(N2262) );
  CMX2X1 U15753 ( .A0(mem_data1[201]), .A1(mem_data1[202]), .S(n3868), .Z(
        n6882) );
  CMXI2X1 U15754 ( .A0(n6882), .A1(n6876), .S(n4065), .Z(n6892) );
  CMX2X1 U15755 ( .A0(n6877), .A1(n6892), .S(n4358), .Z(n6905) );
  CMXI2X1 U15756 ( .A0(n6878), .A1(n6905), .S(n3493), .Z(N2263) );
  CMX2X1 U15757 ( .A0(mem_data1[202]), .A1(mem_data1[203]), .S(n3869), .Z(
        n6888) );
  CMXI2X1 U15758 ( .A0(n6888), .A1(n6879), .S(n4065), .Z(n6895) );
  CMX2X1 U15759 ( .A0(n6880), .A1(n6895), .S(n4358), .Z(n6908) );
  CMXI2X1 U15760 ( .A0(n6881), .A1(n6908), .S(n3493), .Z(N2264) );
  CMX2X1 U15761 ( .A0(mem_data1[203]), .A1(mem_data1[204]), .S(n3870), .Z(
        n6891) );
  CMXI2X1 U15762 ( .A0(n6891), .A1(n6882), .S(n4065), .Z(n6898) );
  CMX2X1 U15763 ( .A0(n6883), .A1(n6898), .S(n4358), .Z(n6911) );
  CMXI2X1 U15764 ( .A0(n6884), .A1(n6911), .S(n3493), .Z(N2265) );
  CMX2X1 U15765 ( .A0(mem_data1[32]), .A1(mem_data1[33]), .S(n3871), .Z(n6956)
         );
  CMXI2X1 U15766 ( .A0(n6956), .A1(n6885), .S(n4065), .Z(n7023) );
  CMX2X1 U15767 ( .A0(n6886), .A1(n7023), .S(n4358), .Z(n7156) );
  CMXI2X1 U15768 ( .A0(n6887), .A1(n7156), .S(n3493), .Z(N2094) );
  CMX2X1 U15769 ( .A0(mem_data1[204]), .A1(mem_data1[205]), .S(n3872), .Z(
        n6894) );
  CMXI2X1 U15770 ( .A0(n6894), .A1(n6888), .S(n4065), .Z(n6901) );
  CMX2X1 U15771 ( .A0(n6889), .A1(n6901), .S(n4358), .Z(n6914) );
  CMXI2X1 U15772 ( .A0(n6890), .A1(n6914), .S(n3493), .Z(N2266) );
  CMX2X1 U15773 ( .A0(mem_data1[205]), .A1(mem_data1[206]), .S(n3873), .Z(
        n6897) );
  CMXI2X1 U15774 ( .A0(n6897), .A1(n6891), .S(n4065), .Z(n6904) );
  CMX2X1 U15775 ( .A0(n6892), .A1(n6904), .S(n4358), .Z(n6917) );
  CMXI2X1 U15776 ( .A0(n6893), .A1(n6917), .S(n3493), .Z(N2267) );
  CMX2X1 U15777 ( .A0(mem_data1[206]), .A1(mem_data1[207]), .S(n3870), .Z(
        n6900) );
  CMXI2X1 U15778 ( .A0(n6900), .A1(n6894), .S(n4064), .Z(n6907) );
  CMX2X1 U15779 ( .A0(n6895), .A1(n6907), .S(n4358), .Z(n6928) );
  CMXI2X1 U15780 ( .A0(n6896), .A1(n6928), .S(n3493), .Z(N2268) );
  CMX2X1 U15781 ( .A0(mem_data1[207]), .A1(mem_data1[208]), .S(n3871), .Z(
        n6903) );
  CMXI2X1 U15782 ( .A0(n6903), .A1(n6897), .S(n4064), .Z(n6910) );
  CMX2X1 U15783 ( .A0(n6898), .A1(n6910), .S(n4358), .Z(n6931) );
  CMXI2X1 U15784 ( .A0(n6899), .A1(n6931), .S(n3493), .Z(N2269) );
  CMX2X1 U15785 ( .A0(mem_data1[208]), .A1(mem_data1[209]), .S(n3874), .Z(
        n6906) );
  CMXI2X1 U15786 ( .A0(n6906), .A1(n6900), .S(n4064), .Z(n6913) );
  CMX2X1 U15787 ( .A0(n6901), .A1(n6913), .S(n4358), .Z(n6934) );
  CMXI2X1 U15788 ( .A0(n6902), .A1(n6934), .S(n3493), .Z(N2270) );
  CMX2X1 U15789 ( .A0(mem_data1[209]), .A1(mem_data1[210]), .S(n3875), .Z(
        n6909) );
  CMXI2X1 U15790 ( .A0(n6909), .A1(n6903), .S(n4064), .Z(n6916) );
  CMX2X1 U15791 ( .A0(n6904), .A1(n6916), .S(n4357), .Z(n6937) );
  CMXI2X1 U15792 ( .A0(n6905), .A1(n6937), .S(n3493), .Z(N2271) );
  CMX2X1 U15793 ( .A0(mem_data1[210]), .A1(mem_data1[211]), .S(n3880), .Z(
        n6912) );
  CMXI2X1 U15794 ( .A0(n6912), .A1(n6906), .S(n4064), .Z(n6927) );
  CMX2X1 U15795 ( .A0(n6907), .A1(n6927), .S(n4357), .Z(n6940) );
  CMXI2X1 U15796 ( .A0(n6908), .A1(n6940), .S(n3492), .Z(N2272) );
  CMX2X1 U15797 ( .A0(mem_data1[211]), .A1(mem_data1[212]), .S(n3881), .Z(
        n6915) );
  CMXI2X1 U15798 ( .A0(n6915), .A1(n6909), .S(n4064), .Z(n6930) );
  CMX2X1 U15799 ( .A0(n6910), .A1(n6930), .S(n4357), .Z(n6943) );
  CMXI2X1 U15800 ( .A0(n6911), .A1(n6943), .S(n3492), .Z(N2273) );
  CMX2X1 U15801 ( .A0(mem_data1[212]), .A1(mem_data1[213]), .S(n3862), .Z(
        n6926) );
  CMXI2X1 U15802 ( .A0(n6926), .A1(n6912), .S(n4064), .Z(n6933) );
  CMX2X1 U15803 ( .A0(n6913), .A1(n6933), .S(n4357), .Z(n6946) );
  CMXI2X1 U15804 ( .A0(n6914), .A1(n6946), .S(n3492), .Z(N2274) );
  CMX2X1 U15805 ( .A0(mem_data1[213]), .A1(mem_data1[214]), .S(n3863), .Z(
        n6929) );
  CMXI2X1 U15806 ( .A0(n6929), .A1(n6915), .S(n4064), .Z(n6936) );
  CMX2X1 U15807 ( .A0(n6916), .A1(n6936), .S(n4357), .Z(n6949) );
  CMXI2X1 U15808 ( .A0(n6917), .A1(n6949), .S(n3495), .Z(N2275) );
  CMX2X1 U15809 ( .A0(mem_data1[33]), .A1(mem_data1[34]), .S(n3873), .Z(n6989)
         );
  CMXI2X1 U15810 ( .A0(n6989), .A1(n6918), .S(n4064), .Z(n7056) );
  CMX2X1 U15811 ( .A0(n6919), .A1(n7056), .S(n4357), .Z(n7189) );
  CMXI2X1 U15812 ( .A0(n6920), .A1(n7189), .S(n3495), .Z(N2095) );
  CMXI2X1 U15813 ( .A0(mem_data1[8]), .A1(mem_data1[7]), .S(n3890), .Z(n7593)
         );
  CMXI2X1 U15814 ( .A0(mem_data1[6]), .A1(mem_data1[5]), .S(n3889), .Z(n7596)
         );
  CMXI2X1 U15815 ( .A0(n7593), .A1(n7596), .S(n4064), .Z(n8265) );
  CMXI2X1 U15816 ( .A0(mem_data1[3]), .A1(mem_data1[4]), .S(n3867), .Z(n7595)
         );
  CMXI2X1 U15817 ( .A0(mem_data1[2]), .A1(mem_data1[1]), .S(n3882), .Z(n6921)
         );
  CMXI2X1 U15818 ( .A0(n7595), .A1(n6921), .S(n4064), .Z(n6922) );
  CMXI2X1 U15819 ( .A0(n8265), .A1(n6922), .S(n3784), .Z(n6925) );
  CMXI2X1 U15820 ( .A0(mem_data1[10]), .A1(mem_data1[9]), .S(n3884), .Z(n7594)
         );
  CMXI2X1 U15821 ( .A0(n6923), .A1(n4430), .S(n4064), .Z(n8264) );
  CMX2X1 U15822 ( .A0(n8264), .A1(n6924), .S(n4357), .Z(n9587) );
  CMXI2X1 U15823 ( .A0(n6925), .A1(n9587), .S(n3495), .Z(N2077) );
  CMX2X1 U15824 ( .A0(mem_data1[214]), .A1(mem_data1[215]), .S(n3874), .Z(
        n6932) );
  CMXI2X1 U15825 ( .A0(n6932), .A1(n6926), .S(n4064), .Z(n6939) );
  CMX2X1 U15826 ( .A0(n6927), .A1(n6939), .S(n4357), .Z(n6952) );
  CMXI2X1 U15827 ( .A0(n6928), .A1(n6952), .S(n3495), .Z(N2276) );
  CMX2X1 U15828 ( .A0(mem_data1[215]), .A1(mem_data1[216]), .S(n3875), .Z(
        n6935) );
  CMXI2X1 U15829 ( .A0(n6935), .A1(n6929), .S(n4064), .Z(n6942) );
  CMX2X1 U15830 ( .A0(n6930), .A1(n6942), .S(n4357), .Z(n6955) );
  CMXI2X1 U15831 ( .A0(n6931), .A1(n6955), .S(n3495), .Z(N2277) );
  CMX2X1 U15832 ( .A0(mem_data1[216]), .A1(mem_data1[217]), .S(n3876), .Z(
        n6938) );
  CMXI2X1 U15833 ( .A0(n6938), .A1(n6932), .S(n4064), .Z(n6945) );
  CMX2X1 U15834 ( .A0(n6933), .A1(n6945), .S(n4357), .Z(n6961) );
  CMXI2X1 U15835 ( .A0(n6934), .A1(n6961), .S(n3495), .Z(N2278) );
  CMX2X1 U15836 ( .A0(mem_data1[217]), .A1(mem_data1[218]), .S(n3876), .Z(
        n6941) );
  CMXI2X1 U15837 ( .A0(n6941), .A1(n6935), .S(n4064), .Z(n6948) );
  CMX2X1 U15838 ( .A0(n6936), .A1(n6948), .S(n4357), .Z(n6964) );
  CMXI2X1 U15839 ( .A0(n6937), .A1(n6964), .S(n3495), .Z(N2279) );
  CMX2X1 U15840 ( .A0(mem_data1[218]), .A1(mem_data1[219]), .S(n3876), .Z(
        n6944) );
  CMXI2X1 U15841 ( .A0(n6944), .A1(n6938), .S(n4063), .Z(n6951) );
  CMX2X1 U15842 ( .A0(n6939), .A1(n6951), .S(n4356), .Z(n6967) );
  CMXI2X1 U15843 ( .A0(n6940), .A1(n6967), .S(n3495), .Z(N2280) );
  CMX2X1 U15844 ( .A0(mem_data1[219]), .A1(mem_data1[220]), .S(n3877), .Z(
        n6947) );
  CMXI2X1 U15845 ( .A0(n6947), .A1(n6941), .S(n4063), .Z(n6954) );
  CMX2X1 U15846 ( .A0(n6942), .A1(n6954), .S(n4356), .Z(n6970) );
  CMXI2X1 U15847 ( .A0(n6943), .A1(n6970), .S(n3495), .Z(N2281) );
  CMX2X1 U15848 ( .A0(mem_data1[220]), .A1(mem_data1[221]), .S(n3878), .Z(
        n6950) );
  CMXI2X1 U15849 ( .A0(n6950), .A1(n6944), .S(n4063), .Z(n6960) );
  CMX2X1 U15850 ( .A0(n6945), .A1(n6960), .S(n4356), .Z(n6973) );
  CMXI2X1 U15851 ( .A0(n6946), .A1(n6973), .S(n3495), .Z(N2282) );
  CMX2X1 U15852 ( .A0(mem_data1[221]), .A1(mem_data1[222]), .S(n3879), .Z(
        n6953) );
  CMXI2X1 U15853 ( .A0(n6953), .A1(n6947), .S(n4063), .Z(n6963) );
  CMX2X1 U15854 ( .A0(n6948), .A1(n6963), .S(n4356), .Z(n6976) );
  CMXI2X1 U15855 ( .A0(n6949), .A1(n6976), .S(n3495), .Z(N2283) );
  CMX2X1 U15856 ( .A0(mem_data1[222]), .A1(mem_data1[223]), .S(n3880), .Z(
        n6959) );
  CMXI2X1 U15857 ( .A0(n6959), .A1(n6950), .S(n4063), .Z(n6966) );
  CMX2X1 U15858 ( .A0(n6951), .A1(n6966), .S(n4356), .Z(n6979) );
  CMXI2X1 U15859 ( .A0(n6952), .A1(n6979), .S(n3494), .Z(N2284) );
  CMX2X1 U15860 ( .A0(mem_data1[223]), .A1(mem_data1[224]), .S(n3881), .Z(
        n6962) );
  CMXI2X1 U15861 ( .A0(n6962), .A1(n6953), .S(n4063), .Z(n6969) );
  CMX2X1 U15862 ( .A0(n6954), .A1(n6969), .S(n4356), .Z(n6982) );
  CMXI2X1 U15863 ( .A0(n6955), .A1(n6982), .S(n3494), .Z(N2285) );
  CMX2X1 U15864 ( .A0(mem_data1[34]), .A1(mem_data1[35]), .S(n3862), .Z(n7022)
         );
  CMXI2X1 U15865 ( .A0(n7022), .A1(n6956), .S(n4063), .Z(n7089) );
  CMX2X1 U15866 ( .A0(n6957), .A1(n7089), .S(n4356), .Z(n7222) );
  CMXI2X1 U15867 ( .A0(n6958), .A1(n7222), .S(n3494), .Z(N2096) );
  CMX2X1 U15868 ( .A0(mem_data1[224]), .A1(mem_data1[225]), .S(n3872), .Z(
        n6965) );
  CMXI2X1 U15869 ( .A0(n6965), .A1(n6959), .S(n4063), .Z(n6972) );
  CMX2X1 U15870 ( .A0(n6960), .A1(n6972), .S(n4356), .Z(n6985) );
  CMXI2X1 U15871 ( .A0(n6961), .A1(n6985), .S(n3494), .Z(N2286) );
  CMX2X1 U15872 ( .A0(mem_data1[225]), .A1(mem_data1[226]), .S(n3873), .Z(
        n6968) );
  CMXI2X1 U15873 ( .A0(n6968), .A1(n6962), .S(n4063), .Z(n6975) );
  CMX2X1 U15874 ( .A0(n6963), .A1(n6975), .S(n4356), .Z(n6988) );
  CMXI2X1 U15875 ( .A0(n6964), .A1(n6988), .S(n3494), .Z(N2287) );
  CMX2X1 U15876 ( .A0(mem_data1[226]), .A1(mem_data1[227]), .S(n3863), .Z(
        n6971) );
  CMXI2X1 U15877 ( .A0(n6971), .A1(n6965), .S(n4063), .Z(n6978) );
  CMX2X1 U15878 ( .A0(n6966), .A1(n6978), .S(n4356), .Z(n6994) );
  CMXI2X1 U15879 ( .A0(n6967), .A1(n6994), .S(n3494), .Z(N2288) );
  CMX2X1 U15880 ( .A0(mem_data1[227]), .A1(mem_data1[228]), .S(n3864), .Z(
        n6974) );
  CMXI2X1 U15881 ( .A0(n6974), .A1(n6968), .S(n4063), .Z(n6981) );
  CMX2X1 U15882 ( .A0(n6969), .A1(n6981), .S(n4356), .Z(n6997) );
  CMXI2X1 U15883 ( .A0(n6970), .A1(n6997), .S(n3494), .Z(N2289) );
  CMX2X1 U15884 ( .A0(mem_data1[228]), .A1(mem_data1[229]), .S(n3864), .Z(
        n6977) );
  CMXI2X1 U15885 ( .A0(n6977), .A1(n6971), .S(n4063), .Z(n6984) );
  CMX2X1 U15886 ( .A0(n6972), .A1(n6984), .S(n4355), .Z(n7000) );
  CMXI2X1 U15887 ( .A0(n6973), .A1(n7000), .S(n3497), .Z(N2290) );
  CMX2X1 U15888 ( .A0(mem_data1[229]), .A1(mem_data1[230]), .S(n3865), .Z(
        n6980) );
  CMXI2X1 U15889 ( .A0(n6980), .A1(n6974), .S(n4063), .Z(n6987) );
  CMX2X1 U15890 ( .A0(n6975), .A1(n6987), .S(n4355), .Z(n7003) );
  CMXI2X1 U15891 ( .A0(n6976), .A1(n7003), .S(n3497), .Z(N2291) );
  CMX2X1 U15892 ( .A0(mem_data1[230]), .A1(mem_data1[231]), .S(n3866), .Z(
        n6983) );
  CMXI2X1 U15893 ( .A0(n6983), .A1(n6977), .S(n4063), .Z(n6993) );
  CMX2X1 U15894 ( .A0(n6978), .A1(n6993), .S(n4355), .Z(n7006) );
  CMXI2X1 U15895 ( .A0(n6979), .A1(n7006), .S(n3497), .Z(N2292) );
  CMX2X1 U15896 ( .A0(mem_data1[231]), .A1(mem_data1[232]), .S(n3867), .Z(
        n6986) );
  CMXI2X1 U15897 ( .A0(n6986), .A1(n6980), .S(n4063), .Z(n6996) );
  CMX2X1 U15898 ( .A0(n6981), .A1(n6996), .S(n4355), .Z(n7009) );
  CMXI2X1 U15899 ( .A0(n6982), .A1(n7009), .S(n3497), .Z(N2293) );
  CMX2X1 U15900 ( .A0(mem_data1[232]), .A1(mem_data1[233]), .S(n3877), .Z(
        n6992) );
  CMXI2X1 U15901 ( .A0(n6992), .A1(n6983), .S(n4063), .Z(n6999) );
  CMX2X1 U15902 ( .A0(n6984), .A1(n6999), .S(n4355), .Z(n7012) );
  CMXI2X1 U15903 ( .A0(n6985), .A1(n7012), .S(n3497), .Z(N2294) );
  CMX2X1 U15904 ( .A0(mem_data1[233]), .A1(mem_data1[234]), .S(n3878), .Z(
        n6995) );
  CMXI2X1 U15905 ( .A0(n6995), .A1(n6986), .S(n4062), .Z(n7002) );
  CMX2X1 U15906 ( .A0(n6987), .A1(n7002), .S(n4355), .Z(n7015) );
  CMXI2X1 U15907 ( .A0(n6988), .A1(n7015), .S(n3497), .Z(N2295) );
  CMX2X1 U15908 ( .A0(mem_data1[35]), .A1(mem_data1[36]), .S(n3879), .Z(n7055)
         );
  CMXI2X1 U15909 ( .A0(n7055), .A1(n6989), .S(n4062), .Z(n7122) );
  CMX2X1 U15910 ( .A0(n6990), .A1(n7122), .S(n4355), .Z(n7255) );
  CMXI2X1 U15911 ( .A0(n6991), .A1(n7255), .S(n3497), .Z(N2097) );
  CMX2X1 U15912 ( .A0(mem_data1[234]), .A1(mem_data1[235]), .S(n3880), .Z(
        n6998) );
  CMXI2X1 U15913 ( .A0(n6998), .A1(n6992), .S(n4062), .Z(n7005) );
  CMX2X1 U15914 ( .A0(n6993), .A1(n7005), .S(n4355), .Z(n7018) );
  CMXI2X1 U15915 ( .A0(n6994), .A1(n7018), .S(n3496), .Z(N2296) );
  CMX2X1 U15916 ( .A0(mem_data1[235]), .A1(mem_data1[236]), .S(n3877), .Z(
        n7001) );
  CMXI2X1 U15917 ( .A0(n7001), .A1(n6995), .S(n4062), .Z(n7008) );
  CMX2X1 U15918 ( .A0(n6996), .A1(n7008), .S(n4355), .Z(n7021) );
  CMXI2X1 U15919 ( .A0(n6997), .A1(n7021), .S(n3496), .Z(N2297) );
  CMX2X1 U15920 ( .A0(mem_data1[236]), .A1(mem_data1[237]), .S(n3865), .Z(
        n7004) );
  CMXI2X1 U15921 ( .A0(n7004), .A1(n6998), .S(n4062), .Z(n7011) );
  CMX2X1 U15922 ( .A0(n6999), .A1(n7011), .S(n4355), .Z(n7027) );
  CMXI2X1 U15923 ( .A0(n7000), .A1(n7027), .S(n3496), .Z(N2298) );
  CMX2X1 U15924 ( .A0(mem_data1[237]), .A1(mem_data1[238]), .S(n3866), .Z(
        n7007) );
  CMXI2X1 U15925 ( .A0(n7007), .A1(n7001), .S(n4062), .Z(n7014) );
  CMX2X1 U15926 ( .A0(n7002), .A1(n7014), .S(n4355), .Z(n7030) );
  CMXI2X1 U15927 ( .A0(n7003), .A1(n7030), .S(n3496), .Z(N2299) );
  CMX2X1 U15928 ( .A0(mem_data1[238]), .A1(mem_data1[239]), .S(n3867), .Z(
        n7010) );
  CMXI2X1 U15929 ( .A0(n7010), .A1(n7004), .S(n4062), .Z(n7017) );
  CMX2X1 U15930 ( .A0(n7005), .A1(n7017), .S(n4354), .Z(n7033) );
  CMXI2X1 U15931 ( .A0(n7006), .A1(n7033), .S(n3496), .Z(N2300) );
  CMX2X1 U15932 ( .A0(mem_data1[239]), .A1(mem_data1[240]), .S(n3868), .Z(
        n7013) );
  CMXI2X1 U15933 ( .A0(n7013), .A1(n7007), .S(n4062), .Z(n7020) );
  CMX2X1 U15934 ( .A0(n7008), .A1(n7020), .S(n4354), .Z(n7036) );
  CMXI2X1 U15935 ( .A0(n7009), .A1(n7036), .S(n3496), .Z(N2301) );
  CMX2X1 U15936 ( .A0(mem_data1[240]), .A1(mem_data1[241]), .S(n3867), .Z(
        n7016) );
  CMXI2X1 U15937 ( .A0(n7016), .A1(n7010), .S(n4062), .Z(n7026) );
  CMX2X1 U15938 ( .A0(n7011), .A1(n7026), .S(n4354), .Z(n7039) );
  CMXI2X1 U15939 ( .A0(n7012), .A1(n7039), .S(n3496), .Z(N2302) );
  CMX2X1 U15940 ( .A0(mem_data1[241]), .A1(mem_data1[242]), .S(n4236), .Z(
        n7019) );
  CMXI2X1 U15941 ( .A0(n7019), .A1(n7013), .S(n4062), .Z(n7029) );
  CMX2X1 U15942 ( .A0(n7014), .A1(n7029), .S(n4354), .Z(n7042) );
  CMXI2X1 U15943 ( .A0(n7015), .A1(n7042), .S(n3496), .Z(N2303) );
  CMX2X1 U15944 ( .A0(mem_data1[242]), .A1(mem_data1[243]), .S(n4236), .Z(
        n7025) );
  CMXI2X1 U15945 ( .A0(n7025), .A1(n7016), .S(n4062), .Z(n7032) );
  CMX2X1 U15946 ( .A0(n7017), .A1(n7032), .S(n4354), .Z(n7045) );
  CMXI2X1 U15947 ( .A0(n7018), .A1(n7045), .S(n3496), .Z(N2304) );
  CMX2X1 U15948 ( .A0(mem_data1[243]), .A1(mem_data1[244]), .S(n4236), .Z(
        n7028) );
  CMXI2X1 U15949 ( .A0(n7028), .A1(n7019), .S(n4062), .Z(n7035) );
  CMX2X1 U15950 ( .A0(n7020), .A1(n7035), .S(n4354), .Z(n7048) );
  CMXI2X1 U15951 ( .A0(n7021), .A1(n7048), .S(n3496), .Z(N2305) );
  CMX2X1 U15952 ( .A0(mem_data1[36]), .A1(mem_data1[37]), .S(n4236), .Z(n7088)
         );
  CMXI2X1 U15953 ( .A0(n7088), .A1(n7022), .S(n4062), .Z(n7155) );
  CMX2X1 U15954 ( .A0(n7023), .A1(n7155), .S(n4354), .Z(n7295) );
  CMXI2X1 U15955 ( .A0(n7024), .A1(n7295), .S(n3496), .Z(N2098) );
  CMX2X1 U15956 ( .A0(mem_data1[244]), .A1(mem_data1[245]), .S(n4236), .Z(
        n7031) );
  CMXI2X1 U15957 ( .A0(n7031), .A1(n7025), .S(n4062), .Z(n7038) );
  CMX2X1 U15958 ( .A0(n7026), .A1(n7038), .S(n4354), .Z(n7051) );
  CMXI2X1 U15959 ( .A0(n7027), .A1(n7051), .S(n3464), .Z(N2306) );
  CMX2X1 U15960 ( .A0(mem_data1[245]), .A1(mem_data1[246]), .S(n4236), .Z(
        n7034) );
  CMXI2X1 U15961 ( .A0(n7034), .A1(n7028), .S(n4062), .Z(n7041) );
  CMX2X1 U15962 ( .A0(n7029), .A1(n7041), .S(n4354), .Z(n7054) );
  CMXI2X1 U15963 ( .A0(n7030), .A1(n7054), .S(n3464), .Z(N2307) );
  CMX2X1 U15964 ( .A0(mem_data1[246]), .A1(mem_data1[247]), .S(n4236), .Z(
        n7037) );
  CMXI2X1 U15965 ( .A0(n7037), .A1(n7031), .S(n4062), .Z(n7044) );
  CMX2X1 U15966 ( .A0(n7032), .A1(n7044), .S(n4354), .Z(n7060) );
  CMXI2X1 U15967 ( .A0(n7033), .A1(n7060), .S(n3464), .Z(N2308) );
  CMX2X1 U15968 ( .A0(mem_data1[247]), .A1(mem_data1[248]), .S(n4236), .Z(
        n7040) );
  CMXI2X1 U15969 ( .A0(n7040), .A1(n7034), .S(n4061), .Z(n7047) );
  CMX2X1 U15970 ( .A0(n7035), .A1(n7047), .S(n4354), .Z(n7063) );
  CMXI2X1 U15971 ( .A0(n7036), .A1(n7063), .S(n3464), .Z(N2309) );
  CMX2X1 U15972 ( .A0(mem_data1[248]), .A1(mem_data1[249]), .S(n4236), .Z(
        n7043) );
  CMXI2X1 U15973 ( .A0(n7043), .A1(n7037), .S(n4061), .Z(n7050) );
  CMX2X1 U15974 ( .A0(n7038), .A1(n7050), .S(n4353), .Z(n7066) );
  CMXI2X1 U15975 ( .A0(n7039), .A1(n7066), .S(n3464), .Z(N2310) );
  CMX2X1 U15976 ( .A0(mem_data1[249]), .A1(mem_data1[250]), .S(n4235), .Z(
        n7046) );
  CMXI2X1 U15977 ( .A0(n7046), .A1(n7040), .S(n4061), .Z(n7053) );
  CMX2X1 U15978 ( .A0(n7041), .A1(n7053), .S(n4353), .Z(n7069) );
  CMXI2X1 U15979 ( .A0(n7042), .A1(n7069), .S(n3464), .Z(N2311) );
  CMX2X1 U15980 ( .A0(mem_data1[250]), .A1(mem_data1[251]), .S(n4235), .Z(
        n7049) );
  CMXI2X1 U15981 ( .A0(n7049), .A1(n7043), .S(n4061), .Z(n7059) );
  CMX2X1 U15982 ( .A0(n7044), .A1(n7059), .S(n4353), .Z(n7072) );
  CMXI2X1 U15983 ( .A0(n7045), .A1(n7072), .S(n3464), .Z(N2312) );
  CMX2X1 U15984 ( .A0(mem_data1[251]), .A1(mem_data1[252]), .S(n4235), .Z(
        n7052) );
  CMXI2X1 U15985 ( .A0(n7052), .A1(n7046), .S(n4061), .Z(n7062) );
  CMX2X1 U15986 ( .A0(n7047), .A1(n7062), .S(n4353), .Z(n7075) );
  CMXI2X1 U15987 ( .A0(n7048), .A1(n7075), .S(n3463), .Z(N2313) );
  CMX2X1 U15988 ( .A0(mem_data1[252]), .A1(mem_data1[253]), .S(n4235), .Z(
        n7058) );
  CMXI2X1 U15989 ( .A0(n7058), .A1(n7049), .S(n4061), .Z(n7065) );
  CMX2X1 U15990 ( .A0(n7050), .A1(n7065), .S(n4362), .Z(n7078) );
  CMXI2X1 U15991 ( .A0(n7051), .A1(n7078), .S(n3463), .Z(N2314) );
  CMX2X1 U15992 ( .A0(mem_data1[253]), .A1(mem_data1[254]), .S(n4235), .Z(
        n7061) );
  CMXI2X1 U15993 ( .A0(n7061), .A1(n7052), .S(n4061), .Z(n7068) );
  CMX2X1 U15994 ( .A0(n7053), .A1(n7068), .S(n3777), .Z(n7081) );
  CMXI2X1 U15995 ( .A0(n7054), .A1(n7081), .S(n3472), .Z(N2315) );
  CMX2X1 U15996 ( .A0(mem_data1[37]), .A1(mem_data1[38]), .S(n4235), .Z(n7121)
         );
  CMXI2X1 U15997 ( .A0(n7121), .A1(n7055), .S(n4061), .Z(n7188) );
  CMX2X1 U15998 ( .A0(n7056), .A1(n7188), .S(n3790), .Z(n7328) );
  CMXI2X1 U15999 ( .A0(n7057), .A1(n7328), .S(n3498), .Z(N2099) );
  CMX2X1 U16000 ( .A0(mem_data1[254]), .A1(mem_data1[255]), .S(n4235), .Z(
        n7064) );
  CMXI2X1 U16001 ( .A0(n7064), .A1(n7058), .S(n4061), .Z(n7071) );
  CMX2X1 U16002 ( .A0(n7059), .A1(n7071), .S(n3791), .Z(n7084) );
  CMXI2X1 U16003 ( .A0(n7060), .A1(n7084), .S(n3498), .Z(N2316) );
  CMX2X1 U16004 ( .A0(mem_data1[255]), .A1(mem_data1[256]), .S(n4235), .Z(
        n7067) );
  CMXI2X1 U16005 ( .A0(n7067), .A1(n7061), .S(n4061), .Z(n7074) );
  CMX2X1 U16006 ( .A0(n7062), .A1(n7074), .S(n3792), .Z(n7087) );
  CMXI2X1 U16007 ( .A0(n7063), .A1(n7087), .S(n3498), .Z(N2317) );
  CMX2X1 U16008 ( .A0(mem_data1[256]), .A1(mem_data1[257]), .S(n4235), .Z(
        n7070) );
  CMXI2X1 U16009 ( .A0(n7070), .A1(n7064), .S(n4061), .Z(n7077) );
  CMX2X1 U16010 ( .A0(n7065), .A1(n7077), .S(n3793), .Z(n7093) );
  CMXI2X1 U16011 ( .A0(n7066), .A1(n7093), .S(n3498), .Z(N2318) );
  CMX2X1 U16012 ( .A0(mem_data1[257]), .A1(mem_data1[258]), .S(n4235), .Z(
        n7073) );
  CMXI2X1 U16013 ( .A0(n7073), .A1(n7067), .S(n4061), .Z(n7080) );
  CMX2X1 U16014 ( .A0(n7068), .A1(n7080), .S(n3794), .Z(n7096) );
  CMXI2X1 U16015 ( .A0(n7069), .A1(n7096), .S(n3497), .Z(N2319) );
  CMX2X1 U16016 ( .A0(mem_data1[258]), .A1(mem_data1[259]), .S(n4235), .Z(
        n7076) );
  CMXI2X1 U16017 ( .A0(n7076), .A1(n7070), .S(n4061), .Z(n7083) );
  CMX2X1 U16018 ( .A0(n7071), .A1(n7083), .S(n3795), .Z(n7099) );
  CMXI2X1 U16019 ( .A0(n7072), .A1(n7099), .S(n3497), .Z(N2320) );
  CMX2X1 U16020 ( .A0(mem_data1[259]), .A1(mem_data1[260]), .S(n4234), .Z(
        n7079) );
  CMXI2X1 U16021 ( .A0(n7079), .A1(n7073), .S(n4061), .Z(n7086) );
  CMX2X1 U16022 ( .A0(n7074), .A1(n7086), .S(n3796), .Z(n7102) );
  CMXI2X1 U16023 ( .A0(n7075), .A1(n7102), .S(n3497), .Z(N2321) );
  CMX2X1 U16024 ( .A0(mem_data1[260]), .A1(mem_data1[261]), .S(n4234), .Z(
        n7082) );
  CMXI2X1 U16025 ( .A0(n7082), .A1(n7076), .S(n4061), .Z(n7092) );
  CMX2X1 U16026 ( .A0(n7077), .A1(n7092), .S(n3797), .Z(n7105) );
  CMXI2X1 U16027 ( .A0(n7078), .A1(n7105), .S(n3497), .Z(N2322) );
  CMX2X1 U16028 ( .A0(mem_data1[261]), .A1(mem_data1[262]), .S(n4234), .Z(
        n7085) );
  CMXI2X1 U16029 ( .A0(n7085), .A1(n7079), .S(n4061), .Z(n7095) );
  CMX2X1 U16030 ( .A0(n7080), .A1(n7095), .S(n3805), .Z(n7108) );
  CMXI2X1 U16031 ( .A0(n7081), .A1(n7108), .S(n3466), .Z(N2323) );
  CMX2X1 U16032 ( .A0(mem_data1[262]), .A1(mem_data1[263]), .S(n4234), .Z(
        n7091) );
  CMXI2X1 U16033 ( .A0(n7091), .A1(n7082), .S(n4060), .Z(n7098) );
  CMX2X1 U16034 ( .A0(n7083), .A1(n7098), .S(n3806), .Z(n7111) );
  CMXI2X1 U16035 ( .A0(n7084), .A1(n7111), .S(n3466), .Z(N2324) );
  CMX2X1 U16036 ( .A0(mem_data1[263]), .A1(mem_data1[264]), .S(n4234), .Z(
        n7094) );
  CMXI2X1 U16037 ( .A0(n7094), .A1(n7085), .S(n4060), .Z(n7101) );
  CMX2X1 U16038 ( .A0(n7086), .A1(n7101), .S(n3808), .Z(n7114) );
  CMXI2X1 U16039 ( .A0(n7087), .A1(n7114), .S(n3466), .Z(N2325) );
  CMX2X1 U16040 ( .A0(mem_data1[38]), .A1(mem_data1[39]), .S(n4234), .Z(n7154)
         );
  CMXI2X1 U16041 ( .A0(n7154), .A1(n7088), .S(n4060), .Z(n7221) );
  CMX2X1 U16042 ( .A0(n7089), .A1(n7221), .S(n3807), .Z(n7361) );
  CMXI2X1 U16043 ( .A0(n7090), .A1(n7361), .S(n3465), .Z(N2100) );
  CMX2X1 U16044 ( .A0(mem_data1[264]), .A1(mem_data1[265]), .S(n4234), .Z(
        n7097) );
  CMXI2X1 U16045 ( .A0(n7097), .A1(n7091), .S(n4060), .Z(n7104) );
  CMX2X1 U16046 ( .A0(n7092), .A1(n7104), .S(n3794), .Z(n7117) );
  CMXI2X1 U16047 ( .A0(n7093), .A1(n7117), .S(n3465), .Z(N2326) );
  CMX2X1 U16048 ( .A0(mem_data1[265]), .A1(mem_data1[266]), .S(n4234), .Z(
        n7100) );
  CMXI2X1 U16049 ( .A0(n7100), .A1(n7094), .S(n4060), .Z(n7107) );
  CMX2X1 U16050 ( .A0(n7095), .A1(n7107), .S(n3795), .Z(n7120) );
  CMXI2X1 U16051 ( .A0(n7096), .A1(n7120), .S(n3465), .Z(N2327) );
  CMX2X1 U16052 ( .A0(mem_data1[266]), .A1(mem_data1[267]), .S(n4234), .Z(
        n7103) );
  CMXI2X1 U16053 ( .A0(n7103), .A1(n7097), .S(n4060), .Z(n7110) );
  CMX2X1 U16054 ( .A0(n7098), .A1(n7110), .S(n3796), .Z(n7126) );
  CMXI2X1 U16055 ( .A0(n7099), .A1(n7126), .S(n3465), .Z(N2328) );
  CMX2X1 U16056 ( .A0(mem_data1[267]), .A1(mem_data1[268]), .S(n4234), .Z(
        n7106) );
  CMXI2X1 U16057 ( .A0(n7106), .A1(n7100), .S(n4060), .Z(n7113) );
  CMX2X1 U16058 ( .A0(n7101), .A1(n7113), .S(n3797), .Z(n7129) );
  CMXI2X1 U16059 ( .A0(n7102), .A1(n7129), .S(n3465), .Z(N2329) );
  CMX2X1 U16060 ( .A0(mem_data1[268]), .A1(mem_data1[269]), .S(n4234), .Z(
        n7109) );
  CMXI2X1 U16061 ( .A0(n7109), .A1(n7103), .S(n4060), .Z(n7116) );
  CMX2X1 U16062 ( .A0(n7104), .A1(n7116), .S(n3805), .Z(n7132) );
  CMXI2X1 U16063 ( .A0(n7105), .A1(n7132), .S(n3465), .Z(N2330) );
  CMX2X1 U16064 ( .A0(mem_data1[269]), .A1(mem_data1[270]), .S(n4233), .Z(
        n7112) );
  CMXI2X1 U16065 ( .A0(n7112), .A1(n7106), .S(n4060), .Z(n7119) );
  CMX2X1 U16066 ( .A0(n7107), .A1(n7119), .S(n3776), .Z(n7135) );
  CMXI2X1 U16067 ( .A0(n7108), .A1(n7135), .S(n3465), .Z(N2331) );
  CMX2X1 U16068 ( .A0(mem_data1[270]), .A1(mem_data1[271]), .S(n4233), .Z(
        n7115) );
  CMXI2X1 U16069 ( .A0(n7115), .A1(n7109), .S(n4060), .Z(n7125) );
  CMX2X1 U16070 ( .A0(n7110), .A1(n7125), .S(n3807), .Z(n7138) );
  CMXI2X1 U16071 ( .A0(n7111), .A1(n7138), .S(n3465), .Z(N2332) );
  CMX2X1 U16072 ( .A0(mem_data1[271]), .A1(mem_data1[272]), .S(n4233), .Z(
        n7118) );
  CMXI2X1 U16073 ( .A0(n7118), .A1(n7112), .S(n4060), .Z(n7128) );
  CMX2X1 U16074 ( .A0(n7113), .A1(n7128), .S(n3808), .Z(n7141) );
  CMXI2X1 U16075 ( .A0(n7114), .A1(n7141), .S(n3307), .Z(N2333) );
  CMX2X1 U16076 ( .A0(mem_data1[272]), .A1(mem_data1[273]), .S(n4233), .Z(
        n7124) );
  CMXI2X1 U16077 ( .A0(n7124), .A1(n7115), .S(n4060), .Z(n7131) );
  CMX2X1 U16078 ( .A0(n7116), .A1(n7131), .S(n3809), .Z(n7144) );
  CMXI2X1 U16079 ( .A0(n7117), .A1(n7144), .S(n3299), .Z(N2334) );
  CMX2X1 U16080 ( .A0(mem_data1[273]), .A1(mem_data1[274]), .S(n4233), .Z(
        n7127) );
  CMXI2X1 U16081 ( .A0(n7127), .A1(n7118), .S(n4060), .Z(n7134) );
  CMX2X1 U16082 ( .A0(n7119), .A1(n7134), .S(n3810), .Z(n7147) );
  CMXI2X1 U16083 ( .A0(n7120), .A1(n7147), .S(n3299), .Z(N2335) );
  CMX2X1 U16084 ( .A0(mem_data1[39]), .A1(mem_data1[40]), .S(n4233), .Z(n7187)
         );
  CMXI2X1 U16085 ( .A0(n7187), .A1(n7121), .S(n4060), .Z(n7254) );
  CMX2X1 U16086 ( .A0(n7122), .A1(n7254), .S(n3811), .Z(n7394) );
  CMXI2X1 U16087 ( .A0(n7123), .A1(n7394), .S(n3299), .Z(N2101) );
  CMX2X1 U16088 ( .A0(mem_data1[274]), .A1(mem_data1[275]), .S(n4233), .Z(
        n7130) );
  CMXI2X1 U16089 ( .A0(n7130), .A1(n7124), .S(n4060), .Z(n7137) );
  CMX2X1 U16090 ( .A0(n7125), .A1(n7137), .S(n3812), .Z(n7150) );
  CMXI2X1 U16091 ( .A0(n7126), .A1(n7150), .S(n3299), .Z(N2336) );
  CMX2X1 U16092 ( .A0(mem_data1[275]), .A1(mem_data1[276]), .S(n4233), .Z(
        n7133) );
  CMXI2X1 U16093 ( .A0(n7133), .A1(n7127), .S(n4060), .Z(n7140) );
  CMX2X1 U16094 ( .A0(n7128), .A1(n7140), .S(n4364), .Z(n7153) );
  CMXI2X1 U16095 ( .A0(n7129), .A1(n7153), .S(n3299), .Z(N2337) );
  CMX2X1 U16096 ( .A0(mem_data1[276]), .A1(mem_data1[277]), .S(n4233), .Z(
        n7136) );
  CMXI2X1 U16097 ( .A0(n7136), .A1(n7130), .S(n4059), .Z(n7143) );
  CMX2X1 U16098 ( .A0(n7131), .A1(n7143), .S(n3771), .Z(n7159) );
  CMXI2X1 U16099 ( .A0(n7132), .A1(n7159), .S(n3299), .Z(N2338) );
  CMX2X1 U16100 ( .A0(mem_data1[277]), .A1(mem_data1[278]), .S(n4233), .Z(
        n7139) );
  CMXI2X1 U16101 ( .A0(n7139), .A1(n7133), .S(n4059), .Z(n7146) );
  CMX2X1 U16102 ( .A0(n7134), .A1(n7146), .S(n3772), .Z(n7162) );
  CMXI2X1 U16103 ( .A0(n7135), .A1(n7162), .S(n3302), .Z(N2339) );
  CMX2X1 U16104 ( .A0(mem_data1[278]), .A1(mem_data1[279]), .S(n4233), .Z(
        n7142) );
  CMXI2X1 U16105 ( .A0(n7142), .A1(n7136), .S(n4059), .Z(n7149) );
  CMX2X1 U16106 ( .A0(n7137), .A1(n7149), .S(n3773), .Z(n7165) );
  CMXI2X1 U16107 ( .A0(n7138), .A1(n7165), .S(n3302), .Z(N2340) );
  CMX2X1 U16108 ( .A0(mem_data1[279]), .A1(mem_data1[280]), .S(n4232), .Z(
        n7145) );
  CMXI2X1 U16109 ( .A0(n7145), .A1(n7139), .S(n4059), .Z(n7152) );
  CMX2X1 U16110 ( .A0(n7140), .A1(n7152), .S(n3774), .Z(n7168) );
  CMXI2X1 U16111 ( .A0(n7141), .A1(n7168), .S(n3302), .Z(N2341) );
  CMX2X1 U16112 ( .A0(mem_data1[280]), .A1(mem_data1[281]), .S(n4232), .Z(
        n7148) );
  CMXI2X1 U16113 ( .A0(n7148), .A1(n7142), .S(n4059), .Z(n7158) );
  CMX2X1 U16114 ( .A0(n7143), .A1(n7158), .S(n3775), .Z(n7171) );
  CMXI2X1 U16115 ( .A0(n7144), .A1(n7171), .S(n3302), .Z(N2342) );
  CMX2X1 U16116 ( .A0(mem_data1[281]), .A1(mem_data1[282]), .S(n4232), .Z(
        n7151) );
  CMXI2X1 U16117 ( .A0(n7151), .A1(n7145), .S(n4059), .Z(n7161) );
  CMX2X1 U16118 ( .A0(n7146), .A1(n7161), .S(n3776), .Z(n7174) );
  CMXI2X1 U16119 ( .A0(n7147), .A1(n7174), .S(n3302), .Z(N2343) );
  CMX2X1 U16120 ( .A0(mem_data1[282]), .A1(mem_data1[283]), .S(n4232), .Z(
        n7157) );
  CMXI2X1 U16121 ( .A0(n7157), .A1(n7148), .S(n4059), .Z(n7164) );
  CMX2X1 U16122 ( .A0(n7149), .A1(n7164), .S(n3777), .Z(n7177) );
  CMXI2X1 U16123 ( .A0(n7150), .A1(n7177), .S(n3302), .Z(N2344) );
  CMX2X1 U16124 ( .A0(mem_data1[283]), .A1(mem_data1[284]), .S(n4232), .Z(
        n7160) );
  CMXI2X1 U16125 ( .A0(n7160), .A1(n7151), .S(n4059), .Z(n7167) );
  CMX2X1 U16126 ( .A0(n7152), .A1(n7167), .S(n3790), .Z(n7180) );
  CMXI2X1 U16127 ( .A0(n7153), .A1(n7180), .S(n3302), .Z(N2345) );
  CMX2X1 U16128 ( .A0(mem_data1[40]), .A1(mem_data1[41]), .S(n4232), .Z(n7220)
         );
  CMXI2X1 U16129 ( .A0(n7220), .A1(n7154), .S(n4059), .Z(n7294) );
  CMX2X1 U16130 ( .A0(n7155), .A1(n7294), .S(n3791), .Z(n7427) );
  CMXI2X1 U16131 ( .A0(n7156), .A1(n7427), .S(n3302), .Z(N2102) );
  CMX2X1 U16132 ( .A0(mem_data1[284]), .A1(mem_data1[285]), .S(n4232), .Z(
        n7163) );
  CMXI2X1 U16133 ( .A0(n7163), .A1(n7157), .S(n4059), .Z(n7170) );
  CMX2X1 U16134 ( .A0(n7158), .A1(n7170), .S(n3809), .Z(n7183) );
  CMXI2X1 U16135 ( .A0(n7159), .A1(n7183), .S(n3301), .Z(N2346) );
  CMX2X1 U16136 ( .A0(mem_data1[285]), .A1(mem_data1[286]), .S(n4232), .Z(
        n7166) );
  CMXI2X1 U16137 ( .A0(n7166), .A1(n7160), .S(n4059), .Z(n7173) );
  CMX2X1 U16138 ( .A0(n7161), .A1(n7173), .S(n3808), .Z(n7186) );
  CMXI2X1 U16139 ( .A0(n7162), .A1(n7186), .S(n3301), .Z(N2347) );
  CMX2X1 U16140 ( .A0(mem_data1[286]), .A1(mem_data1[287]), .S(n4232), .Z(
        n7169) );
  CMXI2X1 U16141 ( .A0(n7169), .A1(n7163), .S(n4059), .Z(n7176) );
  CMX2X1 U16142 ( .A0(n7164), .A1(n7176), .S(n3806), .Z(n7192) );
  CMXI2X1 U16143 ( .A0(n7165), .A1(n7192), .S(n3301), .Z(N2348) );
  CMX2X1 U16144 ( .A0(mem_data1[287]), .A1(mem_data1[288]), .S(n4232), .Z(
        n7172) );
  CMXI2X1 U16145 ( .A0(n7172), .A1(n7166), .S(n4059), .Z(n7179) );
  CMX2X1 U16146 ( .A0(n7167), .A1(n7179), .S(n3807), .Z(n7195) );
  CMXI2X1 U16147 ( .A0(n7168), .A1(n7195), .S(n3301), .Z(N2349) );
  CMX2X1 U16148 ( .A0(mem_data1[288]), .A1(mem_data1[289]), .S(n4232), .Z(
        n7175) );
  CMXI2X1 U16149 ( .A0(n7175), .A1(n7169), .S(n4059), .Z(n7182) );
  CMX2X1 U16150 ( .A0(n7170), .A1(n7182), .S(n3808), .Z(n7198) );
  CMXI2X1 U16151 ( .A0(n7171), .A1(n7198), .S(n3301), .Z(N2350) );
  CMX2X1 U16152 ( .A0(mem_data1[289]), .A1(mem_data1[290]), .S(n4231), .Z(
        n7178) );
  CMXI2X1 U16153 ( .A0(n7178), .A1(n7172), .S(n4059), .Z(n7185) );
  CMX2X1 U16154 ( .A0(n7173), .A1(n7185), .S(n3809), .Z(n7201) );
  CMXI2X1 U16155 ( .A0(n7174), .A1(n7201), .S(n3301), .Z(N2351) );
  CMX2X1 U16156 ( .A0(mem_data1[290]), .A1(mem_data1[291]), .S(n4231), .Z(
        n7181) );
  CMXI2X1 U16157 ( .A0(n7181), .A1(n7175), .S(n4059), .Z(n7191) );
  CMX2X1 U16158 ( .A0(n7176), .A1(n7191), .S(n3810), .Z(n7204) );
  CMXI2X1 U16159 ( .A0(n7177), .A1(n7204), .S(n3301), .Z(N2352) );
  CMX2X1 U16160 ( .A0(mem_data1[291]), .A1(mem_data1[292]), .S(n4231), .Z(
        n7184) );
  CMXI2X1 U16161 ( .A0(n7184), .A1(n7178), .S(n4058), .Z(n7194) );
  CMX2X1 U16162 ( .A0(n7179), .A1(n7194), .S(n3777), .Z(n7207) );
  CMXI2X1 U16163 ( .A0(n7180), .A1(n7207), .S(n3301), .Z(N2353) );
  CMX2X1 U16164 ( .A0(mem_data1[292]), .A1(mem_data1[293]), .S(n4231), .Z(
        n7190) );
  CMXI2X1 U16165 ( .A0(n7190), .A1(n7181), .S(n4058), .Z(n7197) );
  CMX2X1 U16166 ( .A0(n7182), .A1(n7197), .S(n3792), .Z(n7210) );
  CMXI2X1 U16167 ( .A0(n7183), .A1(n7210), .S(n3301), .Z(N2354) );
  CMX2X1 U16168 ( .A0(mem_data1[293]), .A1(mem_data1[294]), .S(n4231), .Z(
        n7193) );
  CMXI2X1 U16169 ( .A0(n7193), .A1(n7184), .S(n4058), .Z(n7200) );
  CMX2X1 U16170 ( .A0(n7185), .A1(n7200), .S(n3793), .Z(n7213) );
  CMXI2X1 U16171 ( .A0(n7186), .A1(n7213), .S(n3301), .Z(N2355) );
  CMX2X1 U16172 ( .A0(mem_data1[41]), .A1(mem_data1[42]), .S(n4231), .Z(n7253)
         );
  CMXI2X1 U16173 ( .A0(n7253), .A1(n7187), .S(n4058), .Z(n7327) );
  CMX2X1 U16174 ( .A0(n7188), .A1(n7327), .S(n3794), .Z(n7460) );
  CMXI2X1 U16175 ( .A0(n7189), .A1(n7460), .S(n3304), .Z(N2103) );
  CMX2X1 U16176 ( .A0(mem_data1[294]), .A1(mem_data1[295]), .S(n4231), .Z(
        n7196) );
  CMXI2X1 U16177 ( .A0(n7196), .A1(n7190), .S(n4058), .Z(n7203) );
  CMX2X1 U16178 ( .A0(n7191), .A1(n7203), .S(n3795), .Z(n7216) );
  CMXI2X1 U16179 ( .A0(n7192), .A1(n7216), .S(n3304), .Z(N2356) );
  CMX2X1 U16180 ( .A0(mem_data1[295]), .A1(mem_data1[296]), .S(n4231), .Z(
        n7199) );
  CMXI2X1 U16181 ( .A0(n7199), .A1(n7193), .S(n4058), .Z(n7206) );
  CMX2X1 U16182 ( .A0(n7194), .A1(n7206), .S(n3796), .Z(n7219) );
  CMXI2X1 U16183 ( .A0(n7195), .A1(n7219), .S(n3304), .Z(N2357) );
  CMX2X1 U16184 ( .A0(mem_data1[296]), .A1(mem_data1[297]), .S(n4231), .Z(
        n7202) );
  CMXI2X1 U16185 ( .A0(n7202), .A1(n7196), .S(n4058), .Z(n7209) );
  CMX2X1 U16186 ( .A0(n7197), .A1(n7209), .S(n3797), .Z(n7225) );
  CMXI2X1 U16187 ( .A0(n7198), .A1(n7225), .S(n3304), .Z(N2358) );
  CMX2X1 U16188 ( .A0(mem_data1[297]), .A1(mem_data1[298]), .S(n4231), .Z(
        n7205) );
  CMXI2X1 U16189 ( .A0(n7205), .A1(n7199), .S(n4058), .Z(n7212) );
  CMX2X1 U16190 ( .A0(n7200), .A1(n7212), .S(n3805), .Z(n7228) );
  CMXI2X1 U16191 ( .A0(n7201), .A1(n7228), .S(n3303), .Z(N2359) );
  CMX2X1 U16192 ( .A0(mem_data1[298]), .A1(mem_data1[299]), .S(n4231), .Z(
        n7208) );
  CMXI2X1 U16193 ( .A0(n7208), .A1(n7202), .S(n4058), .Z(n7215) );
  CMX2X1 U16194 ( .A0(n7203), .A1(n7215), .S(n3806), .Z(n7231) );
  CMXI2X1 U16195 ( .A0(n7204), .A1(n7231), .S(n3303), .Z(N2360) );
  CMX2X1 U16196 ( .A0(mem_data1[299]), .A1(mem_data1[300]), .S(n4230), .Z(
        n7211) );
  CMXI2X1 U16197 ( .A0(n7211), .A1(n7205), .S(n4058), .Z(n7218) );
  CMX2X1 U16198 ( .A0(n7206), .A1(n7218), .S(n3807), .Z(n7234) );
  CMXI2X1 U16199 ( .A0(n7207), .A1(n7234), .S(n3303), .Z(N2361) );
  CMX2X1 U16200 ( .A0(mem_data1[300]), .A1(mem_data1[301]), .S(n4230), .Z(
        n7214) );
  CMXI2X1 U16201 ( .A0(n7214), .A1(n7208), .S(n4058), .Z(n7224) );
  CMX2X1 U16202 ( .A0(n7209), .A1(n7224), .S(n3808), .Z(n7237) );
  CMXI2X1 U16203 ( .A0(n7210), .A1(n7237), .S(n3303), .Z(N2362) );
  CMX2X1 U16204 ( .A0(mem_data1[301]), .A1(mem_data1[302]), .S(n4230), .Z(
        n7217) );
  CMXI2X1 U16205 ( .A0(n7217), .A1(n7211), .S(n4058), .Z(n7227) );
  CMX2X1 U16206 ( .A0(n7212), .A1(n7227), .S(n3809), .Z(n7240) );
  CMXI2X1 U16207 ( .A0(n7213), .A1(n7240), .S(n3303), .Z(N2363) );
  CMX2X1 U16208 ( .A0(mem_data1[302]), .A1(mem_data1[303]), .S(n4230), .Z(
        n7223) );
  CMXI2X1 U16209 ( .A0(n7223), .A1(n7214), .S(n4058), .Z(n7230) );
  CMX2X1 U16210 ( .A0(n7215), .A1(n7230), .S(n3810), .Z(n7243) );
  CMXI2X1 U16211 ( .A0(n7216), .A1(n7243), .S(n3303), .Z(N2364) );
  CMX2X1 U16212 ( .A0(mem_data1[303]), .A1(mem_data1[304]), .S(n4230), .Z(
        n7226) );
  CMXI2X1 U16213 ( .A0(n7226), .A1(n7217), .S(n4058), .Z(n7233) );
  CMX2X1 U16214 ( .A0(n7218), .A1(n7233), .S(n3811), .Z(n7246) );
  CMXI2X1 U16215 ( .A0(n7219), .A1(n7246), .S(n3303), .Z(N2365) );
  CMX2X1 U16216 ( .A0(mem_data1[42]), .A1(mem_data1[43]), .S(n4230), .Z(n7293)
         );
  CMXI2X1 U16217 ( .A0(n7293), .A1(n7220), .S(n4058), .Z(n7360) );
  CMX2X1 U16218 ( .A0(n7221), .A1(n7360), .S(n3812), .Z(n7493) );
  CMXI2X1 U16219 ( .A0(n7222), .A1(n7493), .S(n3303), .Z(N2104) );
  CMX2X1 U16220 ( .A0(mem_data1[304]), .A1(mem_data1[305]), .S(n4230), .Z(
        n7229) );
  CMXI2X1 U16221 ( .A0(n7229), .A1(n7223), .S(n4058), .Z(n7236) );
  CMX2X1 U16222 ( .A0(n7224), .A1(n7236), .S(n4352), .Z(n7249) );
  CMXI2X1 U16223 ( .A0(n7225), .A1(n7249), .S(n3303), .Z(N2366) );
  CMX2X1 U16224 ( .A0(mem_data1[305]), .A1(mem_data1[306]), .S(n4230), .Z(
        n7232) );
  CMXI2X1 U16225 ( .A0(n7232), .A1(n7226), .S(n4057), .Z(n7239) );
  CMX2X1 U16226 ( .A0(n7227), .A1(n7239), .S(n3771), .Z(n7252) );
  CMXI2X1 U16227 ( .A0(n7228), .A1(n7252), .S(n3303), .Z(N2367) );
  CMX2X1 U16228 ( .A0(mem_data1[306]), .A1(mem_data1[307]), .S(n4230), .Z(
        n7235) );
  CMXI2X1 U16229 ( .A0(n7235), .A1(n7229), .S(n4057), .Z(n7242) );
  CMX2X1 U16230 ( .A0(n7230), .A1(n7242), .S(n3810), .Z(n7265) );
  CMXI2X1 U16231 ( .A0(n7231), .A1(n7265), .S(n3303), .Z(N2368) );
  CMX2X1 U16232 ( .A0(mem_data1[307]), .A1(mem_data1[308]), .S(n4230), .Z(
        n7238) );
  CMXI2X1 U16233 ( .A0(n7238), .A1(n7232), .S(n4057), .Z(n7245) );
  CMX2X1 U16234 ( .A0(n7233), .A1(n7245), .S(n3809), .Z(n7268) );
  CMXI2X1 U16235 ( .A0(n7234), .A1(n7268), .S(n3302), .Z(N2369) );
  CMX2X1 U16236 ( .A0(mem_data1[308]), .A1(mem_data1[309]), .S(n4230), .Z(
        n7241) );
  CMXI2X1 U16237 ( .A0(n7241), .A1(n7235), .S(n4057), .Z(n7248) );
  CMX2X1 U16238 ( .A0(n7236), .A1(n7248), .S(n3811), .Z(n7271) );
  CMXI2X1 U16239 ( .A0(n7237), .A1(n7271), .S(n3302), .Z(N2370) );
  CMX2X1 U16240 ( .A0(mem_data1[309]), .A1(mem_data1[310]), .S(n4229), .Z(
        n7244) );
  CMXI2X1 U16241 ( .A0(n7244), .A1(n7238), .S(n4057), .Z(n7251) );
  CMX2X1 U16242 ( .A0(n7239), .A1(n7251), .S(n3812), .Z(n7274) );
  CMXI2X1 U16243 ( .A0(n7240), .A1(n7274), .S(n3302), .Z(N2371) );
  CMX2X1 U16244 ( .A0(mem_data1[310]), .A1(mem_data1[311]), .S(n4229), .Z(
        n7247) );
  CMXI2X1 U16245 ( .A0(n7247), .A1(n7241), .S(n4057), .Z(n7264) );
  CMX2X1 U16246 ( .A0(n7242), .A1(n7264), .S(n4355), .Z(n7277) );
  CMXI2X1 U16247 ( .A0(n7243), .A1(n7277), .S(n3305), .Z(N2372) );
  CMX2X1 U16248 ( .A0(mem_data1[311]), .A1(mem_data1[312]), .S(n4229), .Z(
        n7250) );
  CMXI2X1 U16249 ( .A0(n7250), .A1(n7244), .S(n4057), .Z(n7267) );
  CMX2X1 U16250 ( .A0(n7245), .A1(n7267), .S(n3771), .Z(n7280) );
  CMXI2X1 U16251 ( .A0(n7246), .A1(n7280), .S(n3305), .Z(N2373) );
  CMX2X1 U16252 ( .A0(mem_data1[312]), .A1(mem_data1[313]), .S(n4229), .Z(
        n7263) );
  CMXI2X1 U16253 ( .A0(n7263), .A1(n7247), .S(n4057), .Z(n7270) );
  CMX2X1 U16254 ( .A0(n7248), .A1(n7270), .S(n3772), .Z(n7283) );
  CMXI2X1 U16255 ( .A0(n7249), .A1(n7283), .S(n3305), .Z(N2374) );
  CMX2X1 U16256 ( .A0(mem_data1[313]), .A1(mem_data1[314]), .S(n4229), .Z(
        n7266) );
  CMXI2X1 U16257 ( .A0(n7266), .A1(n7250), .S(n4057), .Z(n7273) );
  CMX2X1 U16258 ( .A0(n7251), .A1(n7273), .S(n3790), .Z(n7286) );
  CMXI2X1 U16259 ( .A0(n7252), .A1(n7286), .S(n3305), .Z(N2375) );
  CMX2X1 U16260 ( .A0(mem_data1[43]), .A1(mem_data1[44]), .S(n4229), .Z(n7326)
         );
  CMXI2X1 U16261 ( .A0(n7326), .A1(n7253), .S(n4057), .Z(n7393) );
  CMX2X1 U16262 ( .A0(n7254), .A1(n7393), .S(n3772), .Z(n7526) );
  CMXI2X1 U16263 ( .A0(n7255), .A1(n7526), .S(n3305), .Z(N2105) );
  CMXI2X1 U16264 ( .A0(n7257), .A1(n7256), .S(n4057), .Z(n8599) );
  CMXI2X1 U16265 ( .A0(n7259), .A1(n7258), .S(n4057), .Z(n7260) );
  CMXI2X1 U16266 ( .A0(n8599), .A1(n7260), .S(n3780), .Z(n7262) );
  CMXI2X1 U16267 ( .A0(n7262), .A1(n7261), .S(n3305), .Z(N2078) );
  CMX2X1 U16268 ( .A0(mem_data1[314]), .A1(mem_data1[315]), .S(n4229), .Z(
        n7269) );
  CMXI2X1 U16269 ( .A0(n7269), .A1(n7263), .S(n4057), .Z(n7276) );
  CMX2X1 U16270 ( .A0(n7264), .A1(n7276), .S(n3773), .Z(n7289) );
  CMXI2X1 U16271 ( .A0(n7265), .A1(n7289), .S(n3305), .Z(N2376) );
  CMX2X1 U16272 ( .A0(mem_data1[315]), .A1(mem_data1[316]), .S(n4229), .Z(
        n7272) );
  CMXI2X1 U16273 ( .A0(n7272), .A1(n7266), .S(n4057), .Z(n7279) );
  CMX2X1 U16274 ( .A0(n7267), .A1(n7279), .S(n3774), .Z(n7292) );
  CMXI2X1 U16275 ( .A0(n7268), .A1(n7292), .S(n3305), .Z(N2377) );
  CMX2X1 U16276 ( .A0(mem_data1[316]), .A1(mem_data1[317]), .S(n4229), .Z(
        n7275) );
  CMXI2X1 U16277 ( .A0(n7275), .A1(n7269), .S(n4057), .Z(n7282) );
  CMX2X1 U16278 ( .A0(n7270), .A1(n7282), .S(n3775), .Z(n7298) );
  CMXI2X1 U16279 ( .A0(n7271), .A1(n7298), .S(n3305), .Z(N2378) );
  CMX2X1 U16280 ( .A0(mem_data1[317]), .A1(mem_data1[318]), .S(n4229), .Z(
        n7278) );
  CMXI2X1 U16281 ( .A0(n7278), .A1(n7272), .S(n4057), .Z(n7285) );
  CMX2X1 U16282 ( .A0(n7273), .A1(n7285), .S(n3776), .Z(n7301) );
  CMXI2X1 U16283 ( .A0(n7274), .A1(n7301), .S(n3305), .Z(N2379) );
  CMX2X1 U16284 ( .A0(mem_data1[318]), .A1(mem_data1[319]), .S(n4229), .Z(
        n7281) );
  CMXI2X1 U16285 ( .A0(n7281), .A1(n7275), .S(n4056), .Z(n7288) );
  CMX2X1 U16286 ( .A0(n7276), .A1(n7288), .S(n3777), .Z(n7304) );
  CMXI2X1 U16287 ( .A0(n7277), .A1(n7304), .S(n3305), .Z(N2380) );
  CMX2X1 U16288 ( .A0(mem_data1[319]), .A1(mem_data1[320]), .S(n4228), .Z(
        n7284) );
  CMXI2X1 U16289 ( .A0(n7284), .A1(n7278), .S(n4056), .Z(n7291) );
  CMX2X1 U16290 ( .A0(n7279), .A1(n7291), .S(n3790), .Z(n7307) );
  CMXI2X1 U16291 ( .A0(n7280), .A1(n7307), .S(n3304), .Z(N2381) );
  CMX2X1 U16292 ( .A0(mem_data1[320]), .A1(mem_data1[321]), .S(n4228), .Z(
        n7287) );
  CMXI2X1 U16293 ( .A0(n7287), .A1(n7281), .S(n4056), .Z(n7297) );
  CMX2X1 U16294 ( .A0(n7282), .A1(n7297), .S(n3791), .Z(n7310) );
  CMXI2X1 U16295 ( .A0(n7283), .A1(n7310), .S(n3304), .Z(N2382) );
  CMX2X1 U16296 ( .A0(mem_data1[321]), .A1(mem_data1[322]), .S(n4228), .Z(
        n7290) );
  CMXI2X1 U16297 ( .A0(n7290), .A1(n7284), .S(n4056), .Z(n7300) );
  CMX2X1 U16298 ( .A0(n7285), .A1(n7300), .S(n3792), .Z(n7313) );
  CMXI2X1 U16299 ( .A0(n7286), .A1(n7313), .S(n3304), .Z(N2383) );
  CMX2X1 U16300 ( .A0(mem_data1[322]), .A1(mem_data1[323]), .S(n4228), .Z(
        n7296) );
  CMXI2X1 U16301 ( .A0(n7296), .A1(n7287), .S(n4056), .Z(n7303) );
  CMX2X1 U16302 ( .A0(n7288), .A1(n7303), .S(n3793), .Z(n7316) );
  CMXI2X1 U16303 ( .A0(n7289), .A1(n7316), .S(n3304), .Z(N2384) );
  CMX2X1 U16304 ( .A0(mem_data1[323]), .A1(mem_data1[324]), .S(n4228), .Z(
        n7299) );
  CMXI2X1 U16305 ( .A0(n7299), .A1(n7290), .S(n4056), .Z(n7306) );
  CMX2X1 U16306 ( .A0(n7291), .A1(n7306), .S(n3794), .Z(n7319) );
  CMXI2X1 U16307 ( .A0(n7292), .A1(n7319), .S(n3304), .Z(N2385) );
  CMX2X1 U16308 ( .A0(mem_data1[44]), .A1(mem_data1[45]), .S(n4228), .Z(n7359)
         );
  CMXI2X1 U16309 ( .A0(n7359), .A1(n7293), .S(n4056), .Z(n7426) );
  CMX2X1 U16310 ( .A0(n7294), .A1(n7426), .S(n3795), .Z(n7559) );
  CMXI2X1 U16311 ( .A0(n7295), .A1(n7559), .S(n3304), .Z(N2106) );
  CMX2X1 U16312 ( .A0(mem_data1[324]), .A1(mem_data1[325]), .S(n4228), .Z(
        n7302) );
  CMXI2X1 U16313 ( .A0(n7302), .A1(n7296), .S(n4056), .Z(n7309) );
  CMX2X1 U16314 ( .A0(n7297), .A1(n7309), .S(n3796), .Z(n7322) );
  CMXI2X1 U16315 ( .A0(n7298), .A1(n7322), .S(n3304), .Z(N2386) );
  CMX2X1 U16316 ( .A0(mem_data1[325]), .A1(mem_data1[326]), .S(n4228), .Z(
        n7305) );
  CMXI2X1 U16317 ( .A0(n7305), .A1(n7299), .S(n4056), .Z(n7312) );
  CMX2X1 U16318 ( .A0(n7300), .A1(n7312), .S(n3797), .Z(n7325) );
  CMXI2X1 U16319 ( .A0(n7301), .A1(n7325), .S(n3307), .Z(N2387) );
  CMX2X1 U16320 ( .A0(mem_data1[326]), .A1(mem_data1[327]), .S(n4228), .Z(
        n7308) );
  CMXI2X1 U16321 ( .A0(n7308), .A1(n7302), .S(n4056), .Z(n7315) );
  CMX2X1 U16322 ( .A0(n7303), .A1(n7315), .S(n3805), .Z(n7331) );
  CMXI2X1 U16323 ( .A0(n7304), .A1(n7331), .S(n3307), .Z(N2388) );
  CMX2X1 U16324 ( .A0(mem_data1[327]), .A1(mem_data1[328]), .S(n4228), .Z(
        n7311) );
  CMXI2X1 U16325 ( .A0(n7311), .A1(n7305), .S(n4056), .Z(n7318) );
  CMX2X1 U16326 ( .A0(n7306), .A1(n7318), .S(n3806), .Z(n7334) );
  CMXI2X1 U16327 ( .A0(n7307), .A1(n7334), .S(n3307), .Z(N2389) );
  CMX2X1 U16328 ( .A0(mem_data1[328]), .A1(mem_data1[329]), .S(n3875), .Z(
        n7314) );
  CMXI2X1 U16329 ( .A0(n7314), .A1(n7308), .S(n4056), .Z(n7321) );
  CMX2X1 U16330 ( .A0(n7309), .A1(n7321), .S(n3811), .Z(n7337) );
  CMXI2X1 U16331 ( .A0(n7310), .A1(n7337), .S(n3307), .Z(N2390) );
  CMX2X1 U16332 ( .A0(mem_data1[329]), .A1(mem_data1[330]), .S(n3869), .Z(
        n7317) );
  CMXI2X1 U16333 ( .A0(n7317), .A1(n7311), .S(n4056), .Z(n7324) );
  CMX2X1 U16334 ( .A0(n7312), .A1(n7324), .S(n3810), .Z(n7340) );
  CMXI2X1 U16335 ( .A0(n7313), .A1(n7340), .S(n3307), .Z(N2391) );
  CMX2X1 U16336 ( .A0(mem_data1[330]), .A1(mem_data1[331]), .S(n3866), .Z(
        n7320) );
  CMXI2X1 U16337 ( .A0(n7320), .A1(n7314), .S(n4056), .Z(n7330) );
  CMX2X1 U16338 ( .A0(n7315), .A1(n7330), .S(n3773), .Z(n7343) );
  CMXI2X1 U16339 ( .A0(n7316), .A1(n7343), .S(n3307), .Z(N2392) );
  CMX2X1 U16340 ( .A0(mem_data1[331]), .A1(mem_data1[332]), .S(n3867), .Z(
        n7323) );
  CMXI2X1 U16341 ( .A0(n7323), .A1(n7317), .S(n4056), .Z(n7333) );
  CMX2X1 U16342 ( .A0(n7318), .A1(n7333), .S(n3774), .Z(n7346) );
  CMXI2X1 U16343 ( .A0(n7319), .A1(n7346), .S(n3307), .Z(N2393) );
  CMX2X1 U16344 ( .A0(mem_data1[332]), .A1(mem_data1[333]), .S(n3868), .Z(
        n7329) );
  CMXI2X1 U16345 ( .A0(n7329), .A1(n7320), .S(n4056), .Z(n7336) );
  CMX2X1 U16346 ( .A0(n7321), .A1(n7336), .S(n3775), .Z(n7349) );
  CMXI2X1 U16347 ( .A0(n7322), .A1(n7349), .S(n3307), .Z(N2394) );
  CMX2X1 U16348 ( .A0(mem_data1[333]), .A1(mem_data1[334]), .S(n3869), .Z(
        n7332) );
  CMXI2X1 U16349 ( .A0(n7332), .A1(n7323), .S(n4055), .Z(n7339) );
  CMX2X1 U16350 ( .A0(n7324), .A1(n7339), .S(n3776), .Z(n7352) );
  CMXI2X1 U16351 ( .A0(n7325), .A1(n7352), .S(n3306), .Z(N2395) );
  CMX2X1 U16352 ( .A0(mem_data1[45]), .A1(mem_data1[46]), .S(n3870), .Z(n7392)
         );
  CMXI2X1 U16353 ( .A0(n7392), .A1(n7326), .S(n4055), .Z(n7459) );
  CMX2X1 U16354 ( .A0(n7327), .A1(n7459), .S(n3811), .Z(n7592) );
  CMXI2X1 U16355 ( .A0(n7328), .A1(n7592), .S(n3306), .Z(N2107) );
  CMX2X1 U16356 ( .A0(mem_data1[334]), .A1(mem_data1[335]), .S(n3871), .Z(
        n7335) );
  CMXI2X1 U16357 ( .A0(n7335), .A1(n7329), .S(n4055), .Z(n7342) );
  CMX2X1 U16358 ( .A0(n7330), .A1(n7342), .S(n3792), .Z(n7355) );
  CMXI2X1 U16359 ( .A0(n7331), .A1(n7355), .S(n3306), .Z(N2396) );
  CMX2X1 U16360 ( .A0(mem_data1[335]), .A1(mem_data1[336]), .S(n3872), .Z(
        n7338) );
  CMXI2X1 U16361 ( .A0(n7338), .A1(n7332), .S(n4055), .Z(n7345) );
  CMX2X1 U16362 ( .A0(n7333), .A1(n7345), .S(n3793), .Z(n7358) );
  CMXI2X1 U16363 ( .A0(n7334), .A1(n7358), .S(n3306), .Z(N2397) );
  CMX2X1 U16364 ( .A0(mem_data1[336]), .A1(mem_data1[337]), .S(n3876), .Z(
        n7341) );
  CMXI2X1 U16365 ( .A0(n7341), .A1(n7335), .S(n4055), .Z(n7348) );
  CMX2X1 U16366 ( .A0(n7336), .A1(n7348), .S(n3794), .Z(n7364) );
  CMXI2X1 U16367 ( .A0(n7337), .A1(n7364), .S(n3306), .Z(N2398) );
  CMX2X1 U16368 ( .A0(mem_data1[337]), .A1(mem_data1[338]), .S(n3877), .Z(
        n7344) );
  CMXI2X1 U16369 ( .A0(n7344), .A1(n7338), .S(n4055), .Z(n7351) );
  CMX2X1 U16370 ( .A0(n7339), .A1(n7351), .S(n3795), .Z(n7367) );
  CMXI2X1 U16371 ( .A0(n7340), .A1(n7367), .S(n3306), .Z(N2399) );
  CMX2X1 U16372 ( .A0(mem_data1[338]), .A1(mem_data1[339]), .S(n3873), .Z(
        n7347) );
  CMXI2X1 U16373 ( .A0(n7347), .A1(n7341), .S(n4055), .Z(n7354) );
  CMX2X1 U16374 ( .A0(n7342), .A1(n7354), .S(n3797), .Z(n7370) );
  CMXI2X1 U16375 ( .A0(n7343), .A1(n7370), .S(n3306), .Z(N2400) );
  CMX2X1 U16376 ( .A0(mem_data1[339]), .A1(mem_data1[340]), .S(n3874), .Z(
        n7350) );
  CMXI2X1 U16377 ( .A0(n7350), .A1(n7344), .S(n4055), .Z(n7357) );
  CMX2X1 U16378 ( .A0(n7345), .A1(n7357), .S(n3805), .Z(n7373) );
  CMXI2X1 U16379 ( .A0(n7346), .A1(n7373), .S(n3306), .Z(N2401) );
  CMX2X1 U16380 ( .A0(mem_data1[340]), .A1(mem_data1[341]), .S(n3876), .Z(
        n7353) );
  CMXI2X1 U16381 ( .A0(n7353), .A1(n7347), .S(n4055), .Z(n7363) );
  CMX2X1 U16382 ( .A0(n7348), .A1(n7363), .S(n3806), .Z(n7376) );
  CMXI2X1 U16383 ( .A0(n7349), .A1(n7376), .S(n3306), .Z(N2402) );
  CMX2X1 U16384 ( .A0(mem_data1[341]), .A1(mem_data1[342]), .S(n3877), .Z(
        n7356) );
  CMXI2X1 U16385 ( .A0(n7356), .A1(n7350), .S(n4055), .Z(n7366) );
  CMX2X1 U16386 ( .A0(n7351), .A1(n7366), .S(n3807), .Z(n7379) );
  CMXI2X1 U16387 ( .A0(n7352), .A1(n7379), .S(n3306), .Z(N2403) );
  CMX2X1 U16388 ( .A0(mem_data1[342]), .A1(mem_data1[343]), .S(n3878), .Z(
        n7362) );
  CMXI2X1 U16389 ( .A0(n7362), .A1(n7353), .S(n4055), .Z(n7369) );
  CMX2X1 U16390 ( .A0(n7354), .A1(n7369), .S(n3808), .Z(n7382) );
  CMXI2X1 U16391 ( .A0(n7355), .A1(n7382), .S(n3309), .Z(N2404) );
  CMX2X1 U16392 ( .A0(mem_data1[343]), .A1(mem_data1[344]), .S(n3879), .Z(
        n7365) );
  CMXI2X1 U16393 ( .A0(n7365), .A1(n7356), .S(n4055), .Z(n7372) );
  CMX2X1 U16394 ( .A0(n7357), .A1(n7372), .S(n3809), .Z(n7385) );
  CMXI2X1 U16395 ( .A0(n7358), .A1(n7385), .S(n3309), .Z(N2405) );
  CMX2X1 U16396 ( .A0(mem_data1[46]), .A1(mem_data1[47]), .S(n3876), .Z(n7425)
         );
  CMXI2X1 U16397 ( .A0(n7425), .A1(n7359), .S(n4055), .Z(n7492) );
  CMX2X1 U16398 ( .A0(n7360), .A1(n7492), .S(n3810), .Z(n7632) );
  CMXI2X1 U16399 ( .A0(n7361), .A1(n7632), .S(n3309), .Z(N2108) );
  CMX2X1 U16400 ( .A0(mem_data1[344]), .A1(mem_data1[345]), .S(n3877), .Z(
        n7368) );
  CMXI2X1 U16401 ( .A0(n7368), .A1(n7362), .S(n4055), .Z(n7375) );
  CMX2X1 U16402 ( .A0(n7363), .A1(n7375), .S(n3811), .Z(n7388) );
  CMXI2X1 U16403 ( .A0(n7364), .A1(n7388), .S(n3309), .Z(N2406) );
  CMX2X1 U16404 ( .A0(mem_data1[345]), .A1(mem_data1[346]), .S(n3878), .Z(
        n7371) );
  CMXI2X1 U16405 ( .A0(n7371), .A1(n7365), .S(n4055), .Z(n7378) );
  CMX2X1 U16406 ( .A0(n7366), .A1(n7378), .S(n3812), .Z(n7391) );
  CMXI2X1 U16407 ( .A0(n7367), .A1(n7391), .S(n3308), .Z(N2407) );
  CMX2X1 U16408 ( .A0(mem_data1[346]), .A1(mem_data1[347]), .S(n3879), .Z(
        n7374) );
  CMXI2X1 U16409 ( .A0(n7374), .A1(n7368), .S(n4055), .Z(n7381) );
  CMX2X1 U16410 ( .A0(n7369), .A1(n7381), .S(n4362), .Z(n7397) );
  CMXI2X1 U16411 ( .A0(n7370), .A1(n7397), .S(n3308), .Z(N2408) );
  CMX2X1 U16412 ( .A0(mem_data1[347]), .A1(mem_data1[348]), .S(n3870), .Z(
        n7377) );
  CMXI2X1 U16413 ( .A0(n7377), .A1(n7371), .S(n4054), .Z(n7384) );
  CMX2X1 U16414 ( .A0(n7372), .A1(n7384), .S(n3771), .Z(n7400) );
  CMXI2X1 U16415 ( .A0(n7373), .A1(n7400), .S(n3308), .Z(N2409) );
  CMX2X1 U16416 ( .A0(mem_data1[348]), .A1(mem_data1[349]), .S(n3873), .Z(
        n7380) );
  CMXI2X1 U16417 ( .A0(n7380), .A1(n7374), .S(n4054), .Z(n7387) );
  CMX2X1 U16418 ( .A0(n7375), .A1(n7387), .S(n3771), .Z(n7403) );
  CMXI2X1 U16419 ( .A0(n7376), .A1(n7403), .S(n3308), .Z(N2410) );
  CMX2X1 U16420 ( .A0(mem_data1[349]), .A1(mem_data1[350]), .S(n3874), .Z(
        n7383) );
  CMXI2X1 U16421 ( .A0(n7383), .A1(n7377), .S(n4054), .Z(n7390) );
  CMX2X1 U16422 ( .A0(n7378), .A1(n7390), .S(n3791), .Z(n7406) );
  CMXI2X1 U16423 ( .A0(n7379), .A1(n7406), .S(n3308), .Z(N2411) );
  CMX2X1 U16424 ( .A0(mem_data1[350]), .A1(mem_data1[351]), .S(n3875), .Z(
        n7386) );
  CMXI2X1 U16425 ( .A0(n7386), .A1(n7380), .S(n4054), .Z(n7396) );
  CMX2X1 U16426 ( .A0(n7381), .A1(n7396), .S(n3805), .Z(n7409) );
  CMXI2X1 U16427 ( .A0(n7382), .A1(n7409), .S(n3308), .Z(N2412) );
  CMX2X1 U16428 ( .A0(mem_data1[351]), .A1(mem_data1[352]), .S(n3876), .Z(
        n7389) );
  CMXI2X1 U16429 ( .A0(n7389), .A1(n7383), .S(n4054), .Z(n7399) );
  CMX2X1 U16430 ( .A0(n7384), .A1(n7399), .S(n3806), .Z(n7412) );
  CMXI2X1 U16431 ( .A0(n7385), .A1(n7412), .S(n3308), .Z(N2413) );
  CMX2X1 U16432 ( .A0(mem_data1[352]), .A1(mem_data1[353]), .S(n3866), .Z(
        n7395) );
  CMXI2X1 U16433 ( .A0(n7395), .A1(n7386), .S(n4054), .Z(n7402) );
  CMX2X1 U16434 ( .A0(n7387), .A1(n7402), .S(n3807), .Z(n7415) );
  CMXI2X1 U16435 ( .A0(n7388), .A1(n7415), .S(n3308), .Z(N2414) );
  CMX2X1 U16436 ( .A0(mem_data1[353]), .A1(mem_data1[354]), .S(n3866), .Z(
        n7398) );
  CMXI2X1 U16437 ( .A0(n7398), .A1(n7389), .S(n4054), .Z(n7405) );
  CMX2X1 U16438 ( .A0(n7390), .A1(n7405), .S(n4375), .Z(n7418) );
  CMXI2X1 U16439 ( .A0(n7391), .A1(n7418), .S(n3308), .Z(N2415) );
  CMX2X1 U16440 ( .A0(mem_data1[47]), .A1(mem_data1[48]), .S(n3867), .Z(n7458)
         );
  CMXI2X1 U16441 ( .A0(n7458), .A1(n7392), .S(n4054), .Z(n7525) );
  CMX2X1 U16442 ( .A0(n7393), .A1(n7525), .S(n4375), .Z(n7665) );
  CMXI2X1 U16443 ( .A0(n7394), .A1(n7665), .S(n3308), .Z(N2109) );
  CMX2X1 U16444 ( .A0(mem_data1[354]), .A1(mem_data1[355]), .S(n3868), .Z(
        n7401) );
  CMXI2X1 U16445 ( .A0(n7401), .A1(n7395), .S(n4054), .Z(n7408) );
  CMX2X1 U16446 ( .A0(n7396), .A1(n7408), .S(n4375), .Z(n7421) );
  CMXI2X1 U16447 ( .A0(n7397), .A1(n7421), .S(n3308), .Z(N2416) );
  CMX2X1 U16448 ( .A0(mem_data1[355]), .A1(mem_data1[356]), .S(n3869), .Z(
        n7404) );
  CMXI2X1 U16449 ( .A0(n7404), .A1(n7398), .S(n4054), .Z(n7411) );
  CMX2X1 U16450 ( .A0(n7399), .A1(n7411), .S(n4375), .Z(n7424) );
  CMXI2X1 U16451 ( .A0(n7400), .A1(n7424), .S(n3307), .Z(N2417) );
  CMX2X1 U16452 ( .A0(mem_data1[356]), .A1(mem_data1[357]), .S(n3870), .Z(
        n7407) );
  CMXI2X1 U16453 ( .A0(n7407), .A1(n7401), .S(n4054), .Z(n7414) );
  CMX2X1 U16454 ( .A0(n7402), .A1(n7414), .S(n4375), .Z(n7430) );
  CMXI2X1 U16455 ( .A0(n7403), .A1(n7430), .S(n3307), .Z(N2418) );
  CMX2X1 U16456 ( .A0(mem_data1[357]), .A1(mem_data1[358]), .S(n3871), .Z(
        n7410) );
  CMXI2X1 U16457 ( .A0(n7410), .A1(n7404), .S(n4054), .Z(n7417) );
  CMX2X1 U16458 ( .A0(n7405), .A1(n7417), .S(n4375), .Z(n7433) );
  CMXI2X1 U16459 ( .A0(n7406), .A1(n7433), .S(n3310), .Z(N2419) );
  CMX2X1 U16460 ( .A0(mem_data1[358]), .A1(mem_data1[359]), .S(n3872), .Z(
        n7413) );
  CMXI2X1 U16461 ( .A0(n7413), .A1(n7407), .S(n4054), .Z(n7420) );
  CMX2X1 U16462 ( .A0(n7408), .A1(n7420), .S(n4375), .Z(n7436) );
  CMXI2X1 U16463 ( .A0(n7409), .A1(n7436), .S(n3310), .Z(N2420) );
  CMX2X1 U16464 ( .A0(mem_data1[359]), .A1(mem_data1[360]), .S(n3872), .Z(
        n7416) );
  CMXI2X1 U16465 ( .A0(n7416), .A1(n7410), .S(n4054), .Z(n7423) );
  CMX2X1 U16466 ( .A0(n7411), .A1(n7423), .S(n4375), .Z(n7439) );
  CMXI2X1 U16467 ( .A0(n7412), .A1(n7439), .S(n3310), .Z(N2421) );
  CMX2X1 U16468 ( .A0(mem_data1[360]), .A1(mem_data1[361]), .S(n3873), .Z(
        n7419) );
  CMXI2X1 U16469 ( .A0(n7419), .A1(n7413), .S(n4054), .Z(n7429) );
  CMX2X1 U16470 ( .A0(n7414), .A1(n7429), .S(n4375), .Z(n7442) );
  CMXI2X1 U16471 ( .A0(n7415), .A1(n7442), .S(n3310), .Z(N2422) );
  CMX2X1 U16472 ( .A0(mem_data1[361]), .A1(mem_data1[362]), .S(n3873), .Z(
        n7422) );
  CMXI2X1 U16473 ( .A0(n7422), .A1(n7416), .S(n4054), .Z(n7432) );
  CMX2X1 U16474 ( .A0(n7417), .A1(n7432), .S(n4375), .Z(n7445) );
  CMXI2X1 U16475 ( .A0(n7418), .A1(n7445), .S(n3310), .Z(N2423) );
  CMX2X1 U16476 ( .A0(mem_data1[362]), .A1(mem_data1[363]), .S(n3874), .Z(
        n7428) );
  CMXI2X1 U16477 ( .A0(n7428), .A1(n7419), .S(n4053), .Z(n7435) );
  CMX2X1 U16478 ( .A0(n7420), .A1(n7435), .S(n4375), .Z(n7448) );
  CMXI2X1 U16479 ( .A0(n7421), .A1(n7448), .S(n3310), .Z(N2424) );
  CMX2X1 U16480 ( .A0(mem_data1[363]), .A1(mem_data1[364]), .S(n3864), .Z(
        n7431) );
  CMXI2X1 U16481 ( .A0(n7431), .A1(n7422), .S(n4053), .Z(n7438) );
  CMX2X1 U16482 ( .A0(n7423), .A1(n7438), .S(n4374), .Z(n7451) );
  CMXI2X1 U16483 ( .A0(n7424), .A1(n7451), .S(n3310), .Z(N2425) );
  CMX2X1 U16484 ( .A0(mem_data1[48]), .A1(mem_data1[49]), .S(n3865), .Z(n7491)
         );
  CMXI2X1 U16485 ( .A0(n7491), .A1(n7425), .S(n4053), .Z(n7558) );
  CMX2X1 U16486 ( .A0(n7426), .A1(n7558), .S(n4374), .Z(n7698) );
  CMXI2X1 U16487 ( .A0(n7427), .A1(n7698), .S(n3310), .Z(N2110) );
  CMX2X1 U16488 ( .A0(mem_data1[364]), .A1(mem_data1[365]), .S(n3866), .Z(
        n7434) );
  CMXI2X1 U16489 ( .A0(n7434), .A1(n7428), .S(n4053), .Z(n7441) );
  CMX2X1 U16490 ( .A0(n7429), .A1(n7441), .S(n4374), .Z(n7454) );
  CMXI2X1 U16491 ( .A0(n7430), .A1(n7454), .S(n3310), .Z(N2426) );
  CMX2X1 U16492 ( .A0(mem_data1[365]), .A1(mem_data1[366]), .S(n3867), .Z(
        n7437) );
  CMXI2X1 U16493 ( .A0(n7437), .A1(n7431), .S(n4053), .Z(n7444) );
  CMX2X1 U16494 ( .A0(n7432), .A1(n7444), .S(n4374), .Z(n7457) );
  CMXI2X1 U16495 ( .A0(n7433), .A1(n7457), .S(n3310), .Z(N2427) );
  CMX2X1 U16496 ( .A0(mem_data1[366]), .A1(mem_data1[367]), .S(n3877), .Z(
        n7440) );
  CMXI2X1 U16497 ( .A0(n7440), .A1(n7434), .S(n4053), .Z(n7447) );
  CMX2X1 U16498 ( .A0(n7435), .A1(n7447), .S(n4374), .Z(n7463) );
  CMXI2X1 U16499 ( .A0(n7436), .A1(n7463), .S(n3310), .Z(N2428) );
  CMX2X1 U16500 ( .A0(mem_data1[367]), .A1(mem_data1[368]), .S(n3878), .Z(
        n7443) );
  CMXI2X1 U16501 ( .A0(n7443), .A1(n7437), .S(n4053), .Z(n7450) );
  CMX2X1 U16502 ( .A0(n7438), .A1(n7450), .S(n4374), .Z(n7466) );
  CMXI2X1 U16503 ( .A0(n7439), .A1(n7466), .S(n3309), .Z(N2429) );
  CMX2X1 U16504 ( .A0(mem_data1[368]), .A1(mem_data1[369]), .S(n3879), .Z(
        n7446) );
  CMXI2X1 U16505 ( .A0(n7446), .A1(n7440), .S(n4053), .Z(n7453) );
  CMX2X1 U16506 ( .A0(n7441), .A1(n7453), .S(n4374), .Z(n7469) );
  CMXI2X1 U16507 ( .A0(n7442), .A1(n7469), .S(n3309), .Z(N2430) );
  CMX2X1 U16508 ( .A0(mem_data1[369]), .A1(mem_data1[370]), .S(n3880), .Z(
        n7449) );
  CMXI2X1 U16509 ( .A0(n7449), .A1(n7443), .S(n4053), .Z(n7456) );
  CMX2X1 U16510 ( .A0(n7444), .A1(n7456), .S(n4374), .Z(n7472) );
  CMXI2X1 U16511 ( .A0(n7445), .A1(n7472), .S(n3309), .Z(N2431) );
  CMX2X1 U16512 ( .A0(mem_data1[370]), .A1(mem_data1[371]), .S(n3867), .Z(
        n7452) );
  CMXI2X1 U16513 ( .A0(n7452), .A1(n7446), .S(n4053), .Z(n7462) );
  CMX2X1 U16514 ( .A0(n7447), .A1(n7462), .S(n4374), .Z(n7475) );
  CMXI2X1 U16515 ( .A0(n7448), .A1(n7475), .S(n3309), .Z(N2432) );
  CMX2X1 U16516 ( .A0(mem_data1[371]), .A1(mem_data1[372]), .S(n3875), .Z(
        n7455) );
  CMXI2X1 U16517 ( .A0(n7455), .A1(n7449), .S(n4053), .Z(n7465) );
  CMX2X1 U16518 ( .A0(n7450), .A1(n7465), .S(n4374), .Z(n7478) );
  CMXI2X1 U16519 ( .A0(n7451), .A1(n7478), .S(n3309), .Z(N2433) );
  CMX2X1 U16520 ( .A0(mem_data1[372]), .A1(mem_data1[373]), .S(n3876), .Z(
        n7461) );
  CMXI2X1 U16521 ( .A0(n7461), .A1(n7452), .S(n4053), .Z(n7468) );
  CMX2X1 U16522 ( .A0(n7453), .A1(n7468), .S(n4374), .Z(n7481) );
  CMXI2X1 U16523 ( .A0(n7454), .A1(n7481), .S(n3309), .Z(N2434) );
  CMX2X1 U16524 ( .A0(mem_data1[373]), .A1(mem_data1[374]), .S(n3877), .Z(
        n7464) );
  CMXI2X1 U16525 ( .A0(n7464), .A1(n7455), .S(n4053), .Z(n7471) );
  CMX2X1 U16526 ( .A0(n7456), .A1(n7471), .S(n4373), .Z(n7484) );
  CMXI2X1 U16527 ( .A0(n7457), .A1(n7484), .S(n3309), .Z(N2435) );
  CMX2X1 U16528 ( .A0(mem_data1[49]), .A1(mem_data1[50]), .S(n3878), .Z(n7524)
         );
  CMXI2X1 U16529 ( .A0(n7524), .A1(n7458), .S(n4053), .Z(n7591) );
  CMX2X1 U16530 ( .A0(n7459), .A1(n7591), .S(n4373), .Z(n7731) );
  CMXI2X1 U16531 ( .A0(n7460), .A1(n7731), .S(n3312), .Z(N2111) );
  CMX2X1 U16532 ( .A0(mem_data1[374]), .A1(mem_data1[375]), .S(n3879), .Z(
        n7467) );
  CMXI2X1 U16533 ( .A0(n7467), .A1(n7461), .S(n4053), .Z(n7474) );
  CMX2X1 U16534 ( .A0(n7462), .A1(n7474), .S(n4373), .Z(n7487) );
  CMXI2X1 U16535 ( .A0(n7463), .A1(n7487), .S(n3312), .Z(N2436) );
  CMX2X1 U16536 ( .A0(mem_data1[375]), .A1(mem_data1[376]), .S(n3880), .Z(
        n7470) );
  CMXI2X1 U16537 ( .A0(n7470), .A1(n7464), .S(n4053), .Z(n7477) );
  CMX2X1 U16538 ( .A0(n7465), .A1(n7477), .S(n4373), .Z(n7490) );
  CMXI2X1 U16539 ( .A0(n7466), .A1(n7490), .S(n3312), .Z(N2437) );
  CMX2X1 U16540 ( .A0(mem_data1[376]), .A1(mem_data1[377]), .S(n3881), .Z(
        n7473) );
  CMXI2X1 U16541 ( .A0(n7473), .A1(n7467), .S(n4052), .Z(n7480) );
  CMX2X1 U16542 ( .A0(n7468), .A1(n7480), .S(n4373), .Z(n7496) );
  CMXI2X1 U16543 ( .A0(n7469), .A1(n7496), .S(n3312), .Z(N2438) );
  CMX2X1 U16544 ( .A0(mem_data1[377]), .A1(mem_data1[378]), .S(n3874), .Z(
        n7476) );
  CMXI2X1 U16545 ( .A0(n7476), .A1(n7470), .S(n4052), .Z(n7483) );
  CMX2X1 U16546 ( .A0(n7471), .A1(n7483), .S(n4373), .Z(n7499) );
  CMXI2X1 U16547 ( .A0(n7472), .A1(n7499), .S(n3312), .Z(N2439) );
  CMX2X1 U16548 ( .A0(mem_data1[378]), .A1(mem_data1[379]), .S(n3875), .Z(
        n7479) );
  CMXI2X1 U16549 ( .A0(n7479), .A1(n7473), .S(n4052), .Z(n7486) );
  CMX2X1 U16550 ( .A0(n7474), .A1(n7486), .S(n4373), .Z(n7502) );
  CMXI2X1 U16551 ( .A0(n7475), .A1(n7502), .S(n3312), .Z(N2440) );
  CMX2X1 U16552 ( .A0(mem_data1[379]), .A1(mem_data1[380]), .S(n3862), .Z(
        n7482) );
  CMXI2X1 U16553 ( .A0(n7482), .A1(n7476), .S(n4052), .Z(n7489) );
  CMX2X1 U16554 ( .A0(n7477), .A1(n7489), .S(n4373), .Z(n7505) );
  CMXI2X1 U16555 ( .A0(n7478), .A1(n7505), .S(n3312), .Z(N2441) );
  CMX2X1 U16556 ( .A0(mem_data1[380]), .A1(mem_data1[381]), .S(n3863), .Z(
        n7485) );
  CMXI2X1 U16557 ( .A0(n7485), .A1(n7479), .S(n4052), .Z(n7495) );
  CMX2X1 U16558 ( .A0(n7480), .A1(n7495), .S(n4373), .Z(n7508) );
  CMXI2X1 U16559 ( .A0(n7481), .A1(n7508), .S(n3311), .Z(N2442) );
  CMX2X1 U16560 ( .A0(mem_data1[381]), .A1(mem_data1[382]), .S(n3868), .Z(
        n7488) );
  CMXI2X1 U16561 ( .A0(n7488), .A1(n7482), .S(n4052), .Z(n7498) );
  CMX2X1 U16562 ( .A0(n7483), .A1(n7498), .S(n4373), .Z(n7511) );
  CMXI2X1 U16563 ( .A0(n7484), .A1(n7511), .S(n3311), .Z(N2443) );
  CMX2X1 U16564 ( .A0(mem_data1[382]), .A1(mem_data1[383]), .S(n3869), .Z(
        n7494) );
  CMXI2X1 U16565 ( .A0(n7494), .A1(n7485), .S(n4052), .Z(n7501) );
  CMX2X1 U16566 ( .A0(n7486), .A1(n7501), .S(n4373), .Z(n7514) );
  CMXI2X1 U16567 ( .A0(n7487), .A1(n7514), .S(n3311), .Z(N2444) );
  CMX2X1 U16568 ( .A0(mem_data1[383]), .A1(mem_data1[384]), .S(n3870), .Z(
        n7497) );
  CMXI2X1 U16569 ( .A0(n7497), .A1(n7488), .S(n4052), .Z(n7504) );
  CMX2X1 U16570 ( .A0(n7489), .A1(n7504), .S(n4372), .Z(n7517) );
  CMXI2X1 U16571 ( .A0(n7490), .A1(n7517), .S(n3311), .Z(N2445) );
  CMX2X1 U16572 ( .A0(mem_data1[50]), .A1(mem_data1[51]), .S(n3871), .Z(n7557)
         );
  CMXI2X1 U16573 ( .A0(n7557), .A1(n7491), .S(n4052), .Z(n7631) );
  CMX2X1 U16574 ( .A0(n7492), .A1(n7631), .S(n4372), .Z(n7764) );
  CMXI2X1 U16575 ( .A0(n7493), .A1(n7764), .S(n3311), .Z(N2112) );
  CMX2X1 U16576 ( .A0(mem_data1[384]), .A1(mem_data1[385]), .S(n3881), .Z(
        n7500) );
  CMXI2X1 U16577 ( .A0(n7500), .A1(n7494), .S(n4052), .Z(n7507) );
  CMX2X1 U16578 ( .A0(n7495), .A1(n7507), .S(n4372), .Z(n7520) );
  CMXI2X1 U16579 ( .A0(n7496), .A1(n7520), .S(n3311), .Z(N2446) );
  CMX2X1 U16580 ( .A0(mem_data1[385]), .A1(mem_data1[386]), .S(n3862), .Z(
        n7503) );
  CMXI2X1 U16581 ( .A0(n7503), .A1(n7497), .S(n4052), .Z(n7510) );
  CMX2X1 U16582 ( .A0(n7498), .A1(n7510), .S(n4372), .Z(n7523) );
  CMXI2X1 U16583 ( .A0(n7499), .A1(n7523), .S(n3311), .Z(N2447) );
  CMX2X1 U16584 ( .A0(mem_data1[386]), .A1(mem_data1[387]), .S(n3863), .Z(
        n7506) );
  CMXI2X1 U16585 ( .A0(n7506), .A1(n7500), .S(n4052), .Z(n7513) );
  CMX2X1 U16586 ( .A0(n7501), .A1(n7513), .S(n4372), .Z(n7529) );
  CMXI2X1 U16587 ( .A0(n7502), .A1(n7529), .S(n3311), .Z(N2448) );
  CMX2X1 U16588 ( .A0(mem_data1[387]), .A1(mem_data1[388]), .S(n3864), .Z(
        n7509) );
  CMXI2X1 U16589 ( .A0(n7509), .A1(n7503), .S(n4052), .Z(n7516) );
  CMX2X1 U16590 ( .A0(n7504), .A1(n7516), .S(n4372), .Z(n7532) );
  CMXI2X1 U16591 ( .A0(n7505), .A1(n7532), .S(n3311), .Z(N2449) );
  CMX2X1 U16592 ( .A0(mem_data1[388]), .A1(mem_data1[389]), .S(n3868), .Z(
        n7512) );
  CMXI2X1 U16593 ( .A0(n7512), .A1(n7506), .S(n4052), .Z(n7519) );
  CMX2X1 U16594 ( .A0(n7507), .A1(n7519), .S(n4372), .Z(n7535) );
  CMXI2X1 U16595 ( .A0(n7508), .A1(n7535), .S(n3311), .Z(N2450) );
  CMX2X1 U16596 ( .A0(mem_data1[389]), .A1(mem_data1[390]), .S(n3864), .Z(
        n7515) );
  CMXI2X1 U16597 ( .A0(n7515), .A1(n7509), .S(n4052), .Z(n7522) );
  CMX2X1 U16598 ( .A0(n7510), .A1(n7522), .S(n4372), .Z(n7538) );
  CMXI2X1 U16599 ( .A0(n7511), .A1(n7538), .S(n3311), .Z(N2451) );
  CMX2X1 U16600 ( .A0(mem_data1[390]), .A1(mem_data1[391]), .S(n3865), .Z(
        n7518) );
  CMXI2X1 U16601 ( .A0(n7518), .A1(n7512), .S(n4052), .Z(n7528) );
  CMX2X1 U16602 ( .A0(n7513), .A1(n7528), .S(n4372), .Z(n7541) );
  CMXI2X1 U16603 ( .A0(n7514), .A1(n7541), .S(n3314), .Z(N2452) );
  CMX2X1 U16604 ( .A0(mem_data1[391]), .A1(mem_data1[392]), .S(n3866), .Z(
        n7521) );
  CMXI2X1 U16605 ( .A0(n7521), .A1(n7515), .S(n4051), .Z(n7531) );
  CMX2X1 U16606 ( .A0(n7516), .A1(n7531), .S(n4372), .Z(n7544) );
  CMXI2X1 U16607 ( .A0(n7517), .A1(n7544), .S(n3314), .Z(N2453) );
  CMX2X1 U16608 ( .A0(mem_data1[392]), .A1(mem_data1[393]), .S(n3867), .Z(
        n7527) );
  CMXI2X1 U16609 ( .A0(n7527), .A1(n7518), .S(n4051), .Z(n7534) );
  CMX2X1 U16610 ( .A0(n7519), .A1(n7534), .S(n4372), .Z(n7547) );
  CMXI2X1 U16611 ( .A0(n7520), .A1(n7547), .S(n3314), .Z(N2454) );
  CMX2X1 U16612 ( .A0(mem_data1[393]), .A1(mem_data1[394]), .S(n3868), .Z(
        n7530) );
  CMXI2X1 U16613 ( .A0(n7530), .A1(n7521), .S(n4051), .Z(n7537) );
  CMX2X1 U16614 ( .A0(n7522), .A1(n7537), .S(n4371), .Z(n7550) );
  CMXI2X1 U16615 ( .A0(n7523), .A1(n7550), .S(n3313), .Z(N2455) );
  CMX2X1 U16616 ( .A0(mem_data1[51]), .A1(mem_data1[52]), .S(n3869), .Z(n7590)
         );
  CMXI2X1 U16617 ( .A0(n7590), .A1(n7524), .S(n4051), .Z(n7664) );
  CMX2X1 U16618 ( .A0(n7525), .A1(n7664), .S(n4371), .Z(n7797) );
  CMXI2X1 U16619 ( .A0(n7526), .A1(n7797), .S(n3313), .Z(N2113) );
  CMX2X1 U16620 ( .A0(mem_data1[394]), .A1(mem_data1[395]), .S(n3870), .Z(
        n7533) );
  CMXI2X1 U16621 ( .A0(n7533), .A1(n7527), .S(n4051), .Z(n7540) );
  CMX2X1 U16622 ( .A0(n7528), .A1(n7540), .S(n4371), .Z(n7553) );
  CMXI2X1 U16623 ( .A0(n7529), .A1(n7553), .S(n3313), .Z(N2456) );
  CMX2X1 U16624 ( .A0(mem_data1[395]), .A1(mem_data1[396]), .S(n3876), .Z(
        n7536) );
  CMXI2X1 U16625 ( .A0(n7536), .A1(n7530), .S(n4051), .Z(n7543) );
  CMX2X1 U16626 ( .A0(n7531), .A1(n7543), .S(n4371), .Z(n7556) );
  CMXI2X1 U16627 ( .A0(n7532), .A1(n7556), .S(n3313), .Z(N2457) );
  CMX2X1 U16628 ( .A0(mem_data1[396]), .A1(mem_data1[397]), .S(n3877), .Z(
        n7539) );
  CMXI2X1 U16629 ( .A0(n7539), .A1(n7533), .S(n4051), .Z(n7546) );
  CMX2X1 U16630 ( .A0(n7534), .A1(n7546), .S(n4371), .Z(n7562) );
  CMXI2X1 U16631 ( .A0(n7535), .A1(n7562), .S(n3313), .Z(N2458) );
  CMX2X1 U16632 ( .A0(mem_data1[397]), .A1(mem_data1[398]), .S(n3871), .Z(
        n7542) );
  CMXI2X1 U16633 ( .A0(n7542), .A1(n7536), .S(n4051), .Z(n7549) );
  CMX2X1 U16634 ( .A0(n7537), .A1(n7549), .S(n4371), .Z(n7565) );
  CMXI2X1 U16635 ( .A0(n7538), .A1(n7565), .S(n3313), .Z(N2459) );
  CMX2X1 U16636 ( .A0(mem_data1[398]), .A1(mem_data1[399]), .S(n3872), .Z(
        n7545) );
  CMXI2X1 U16637 ( .A0(n7545), .A1(n7539), .S(n4051), .Z(n7552) );
  CMX2X1 U16638 ( .A0(n7540), .A1(n7552), .S(n4371), .Z(n7568) );
  CMXI2X1 U16639 ( .A0(n7541), .A1(n7568), .S(n3313), .Z(N2460) );
  CMX2X1 U16640 ( .A0(mem_data1[399]), .A1(mem_data1[400]), .S(n3872), .Z(
        n7548) );
  CMXI2X1 U16641 ( .A0(n7548), .A1(n7542), .S(n4051), .Z(n7555) );
  CMX2X1 U16642 ( .A0(n7543), .A1(n7555), .S(n4371), .Z(n7571) );
  CMXI2X1 U16643 ( .A0(n7544), .A1(n7571), .S(n3313), .Z(N2461) );
  CMX2X1 U16644 ( .A0(mem_data1[400]), .A1(mem_data1[401]), .S(n3873), .Z(
        n7551) );
  CMXI2X1 U16645 ( .A0(n7551), .A1(n7545), .S(n4051), .Z(n7561) );
  CMX2X1 U16646 ( .A0(n7546), .A1(n7561), .S(n4371), .Z(n7574) );
  CMXI2X1 U16647 ( .A0(n7547), .A1(n7574), .S(n3313), .Z(N2462) );
  CMX2X1 U16648 ( .A0(mem_data1[401]), .A1(mem_data1[402]), .S(n3874), .Z(
        n7554) );
  CMXI2X1 U16649 ( .A0(n7554), .A1(n7548), .S(n4051), .Z(n7564) );
  CMX2X1 U16650 ( .A0(n7549), .A1(n7564), .S(n4371), .Z(n7577) );
  CMXI2X1 U16651 ( .A0(n7550), .A1(n7577), .S(n3313), .Z(N2463) );
  CMX2X1 U16652 ( .A0(mem_data1[402]), .A1(mem_data1[403]), .S(n3875), .Z(
        n7560) );
  CMXI2X1 U16653 ( .A0(n7560), .A1(n7551), .S(n4051), .Z(n7567) );
  CMX2X1 U16654 ( .A0(n7552), .A1(n7567), .S(n4371), .Z(n7580) );
  CMXI2X1 U16655 ( .A0(n7553), .A1(n7580), .S(n3313), .Z(N2464) );
  CMX2X1 U16656 ( .A0(mem_data1[403]), .A1(mem_data1[404]), .S(n3865), .Z(
        n7563) );
  CMXI2X1 U16657 ( .A0(n7563), .A1(n7554), .S(n4051), .Z(n7570) );
  CMX2X1 U16658 ( .A0(n7555), .A1(n7570), .S(n4370), .Z(n7583) );
  CMXI2X1 U16659 ( .A0(n7556), .A1(n7583), .S(n3312), .Z(N2465) );
  CMX2X1 U16660 ( .A0(mem_data1[52]), .A1(mem_data1[53]), .S(n3866), .Z(n7630)
         );
  CMXI2X1 U16661 ( .A0(n7630), .A1(n7557), .S(n4051), .Z(n7697) );
  CMX2X1 U16662 ( .A0(n7558), .A1(n7697), .S(n4370), .Z(n7830) );
  CMXI2X1 U16663 ( .A0(n7559), .A1(n7830), .S(n3312), .Z(N2114) );
  CMX2X1 U16664 ( .A0(mem_data1[404]), .A1(mem_data1[405]), .S(n3867), .Z(
        n7566) );
  CMXI2X1 U16665 ( .A0(n7566), .A1(n7560), .S(n4051), .Z(n7573) );
  CMX2X1 U16666 ( .A0(n7561), .A1(n7573), .S(n4370), .Z(n7586) );
  CMXI2X1 U16667 ( .A0(n7562), .A1(n7586), .S(n3312), .Z(N2466) );
  CMX2X1 U16668 ( .A0(mem_data1[405]), .A1(mem_data1[406]), .S(n3868), .Z(
        n7569) );
  CMXI2X1 U16669 ( .A0(n7569), .A1(n7563), .S(n4050), .Z(n7576) );
  CMX2X1 U16670 ( .A0(n7564), .A1(n7576), .S(n4370), .Z(n7589) );
  CMXI2X1 U16671 ( .A0(n7565), .A1(n7589), .S(n3312), .Z(N2467) );
  CMX2X1 U16672 ( .A0(mem_data1[406]), .A1(mem_data1[407]), .S(n3869), .Z(
        n7572) );
  CMXI2X1 U16673 ( .A0(n7572), .A1(n7566), .S(n4050), .Z(n7579) );
  CMX2X1 U16674 ( .A0(n7567), .A1(n7579), .S(n4370), .Z(n7602) );
  CMXI2X1 U16675 ( .A0(n7568), .A1(n7602), .S(n3481), .Z(N2468) );
  CMX2X1 U16676 ( .A0(mem_data1[407]), .A1(mem_data1[408]), .S(n3873), .Z(
        n7575) );
  CMXI2X1 U16677 ( .A0(n7575), .A1(n7569), .S(n4050), .Z(n7582) );
  CMX2X1 U16678 ( .A0(n7570), .A1(n7582), .S(n4370), .Z(n7605) );
  CMXI2X1 U16679 ( .A0(n7571), .A1(n7605), .S(n3489), .Z(N2469) );
  CMX2X1 U16680 ( .A0(mem_data1[408]), .A1(mem_data1[409]), .S(n3874), .Z(
        n7578) );
  CMXI2X1 U16681 ( .A0(n7578), .A1(n7572), .S(n4050), .Z(n7585) );
  CMX2X1 U16682 ( .A0(n7573), .A1(n7585), .S(n4370), .Z(n7608) );
  CMXI2X1 U16683 ( .A0(n7574), .A1(n7608), .S(n3498), .Z(N2470) );
  CMX2X1 U16684 ( .A0(mem_data1[409]), .A1(mem_data1[410]), .S(n3875), .Z(
        n7581) );
  CMXI2X1 U16685 ( .A0(n7581), .A1(n7575), .S(n4050), .Z(n7588) );
  CMX2X1 U16686 ( .A0(n7576), .A1(n7588), .S(n4370), .Z(n7611) );
  CMXI2X1 U16687 ( .A0(n7577), .A1(n7611), .S(n3332), .Z(N2471) );
  CMX2X1 U16688 ( .A0(mem_data1[410]), .A1(mem_data1[411]), .S(n3876), .Z(
        n7584) );
  CMXI2X1 U16689 ( .A0(n7584), .A1(n7578), .S(n4050), .Z(n7601) );
  CMX2X1 U16690 ( .A0(n7579), .A1(n7601), .S(n4370), .Z(n7614) );
  CMXI2X1 U16691 ( .A0(n7580), .A1(n7614), .S(n3315), .Z(N2472) );
  CMX2X1 U16692 ( .A0(mem_data1[411]), .A1(mem_data1[412]), .S(n3877), .Z(
        n7587) );
  CMXI2X1 U16693 ( .A0(n7587), .A1(n7581), .S(n4050), .Z(n7604) );
  CMX2X1 U16694 ( .A0(n7582), .A1(n7604), .S(n4370), .Z(n7617) );
  CMXI2X1 U16695 ( .A0(n7583), .A1(n7617), .S(n3315), .Z(N2473) );
  CMX2X1 U16696 ( .A0(mem_data1[412]), .A1(mem_data1[413]), .S(n4236), .Z(
        n7600) );
  CMXI2X1 U16697 ( .A0(n7600), .A1(n7584), .S(n4050), .Z(n7607) );
  CMX2X1 U16698 ( .A0(n7585), .A1(n7607), .S(n4370), .Z(n7620) );
  CMXI2X1 U16699 ( .A0(n7586), .A1(n7620), .S(n3315), .Z(N2474) );
  CMX2X1 U16700 ( .A0(mem_data1[413]), .A1(mem_data1[414]), .S(n4228), .Z(
        n7603) );
  CMXI2X1 U16701 ( .A0(n7603), .A1(n7587), .S(n4050), .Z(n7610) );
  CMX2X1 U16702 ( .A0(n7588), .A1(n7610), .S(n4369), .Z(n7623) );
  CMXI2X1 U16703 ( .A0(n7589), .A1(n7623), .S(n3315), .Z(N2475) );
  CMX2X1 U16704 ( .A0(mem_data1[53]), .A1(mem_data1[54]), .S(n3876), .Z(n7663)
         );
  CMXI2X1 U16705 ( .A0(n7663), .A1(n7590), .S(n4050), .Z(n7730) );
  CMX2X1 U16706 ( .A0(n7591), .A1(n7730), .S(n4369), .Z(n7863) );
  CMXI2X1 U16707 ( .A0(n7592), .A1(n7863), .S(n3315), .Z(N2115) );
  CMXI2X1 U16708 ( .A0(n7594), .A1(n7593), .S(n4050), .Z(n8933) );
  CMXI2X1 U16709 ( .A0(n7596), .A1(n7595), .S(n4050), .Z(n7597) );
  CMXI2X1 U16710 ( .A0(n8933), .A1(n7597), .S(n3785), .Z(n7599) );
  CMXI2X1 U16711 ( .A0(n7599), .A1(n7598), .S(n3315), .Z(N2079) );
  CMX2X1 U16712 ( .A0(mem_data1[414]), .A1(mem_data1[415]), .S(n3876), .Z(
        n7606) );
  CMXI2X1 U16713 ( .A0(n7606), .A1(n7600), .S(n4050), .Z(n7613) );
  CMX2X1 U16714 ( .A0(n7601), .A1(n7613), .S(n4369), .Z(n7626) );
  CMXI2X1 U16715 ( .A0(n7602), .A1(n7626), .S(n3314), .Z(N2476) );
  CMX2X1 U16716 ( .A0(mem_data1[415]), .A1(mem_data1[416]), .S(n3877), .Z(
        n7609) );
  CMXI2X1 U16717 ( .A0(n7609), .A1(n7603), .S(n4050), .Z(n7616) );
  CMX2X1 U16718 ( .A0(n7604), .A1(n7616), .S(n4369), .Z(n7629) );
  CMXI2X1 U16719 ( .A0(n7605), .A1(n7629), .S(n3314), .Z(N2477) );
  CMX2X1 U16720 ( .A0(mem_data1[416]), .A1(mem_data1[417]), .S(n3878), .Z(
        n7612) );
  CMXI2X1 U16721 ( .A0(n7612), .A1(n7606), .S(n4050), .Z(n7619) );
  CMX2X1 U16722 ( .A0(n7607), .A1(n7619), .S(n4369), .Z(n7635) );
  CMXI2X1 U16723 ( .A0(n7608), .A1(n7635), .S(n3314), .Z(N2478) );
  CMX2X1 U16724 ( .A0(mem_data1[417]), .A1(mem_data1[418]), .S(n3879), .Z(
        n7615) );
  CMXI2X1 U16725 ( .A0(n7615), .A1(n7609), .S(n4050), .Z(n7622) );
  CMX2X1 U16726 ( .A0(n7610), .A1(n7622), .S(n4369), .Z(n7638) );
  CMXI2X1 U16727 ( .A0(n7611), .A1(n7638), .S(n3314), .Z(N2479) );
  CMX2X1 U16728 ( .A0(mem_data1[418]), .A1(mem_data1[419]), .S(n3869), .Z(
        n7618) );
  CMXI2X1 U16729 ( .A0(n7618), .A1(n7612), .S(n4049), .Z(n7625) );
  CMX2X1 U16730 ( .A0(n7613), .A1(n7625), .S(n4369), .Z(n7641) );
  CMXI2X1 U16731 ( .A0(n7614), .A1(n7641), .S(n3314), .Z(N2480) );
  CMX2X1 U16732 ( .A0(mem_data1[419]), .A1(mem_data1[420]), .S(n3870), .Z(
        n7621) );
  CMXI2X1 U16733 ( .A0(n7621), .A1(n7615), .S(n4049), .Z(n7628) );
  CMX2X1 U16734 ( .A0(n7616), .A1(n7628), .S(n4369), .Z(n7644) );
  CMXI2X1 U16735 ( .A0(n7617), .A1(n7644), .S(n3314), .Z(N2481) );
  CMX2X1 U16736 ( .A0(mem_data1[420]), .A1(mem_data1[421]), .S(n3871), .Z(
        n7624) );
  CMXI2X1 U16737 ( .A0(n7624), .A1(n7618), .S(n4049), .Z(n7634) );
  CMX2X1 U16738 ( .A0(n7619), .A1(n7634), .S(n4369), .Z(n7647) );
  CMXI2X1 U16739 ( .A0(n7620), .A1(n7647), .S(n3314), .Z(N2482) );
  CMX2X1 U16740 ( .A0(mem_data1[421]), .A1(mem_data1[422]), .S(n3872), .Z(
        n7627) );
  CMXI2X1 U16741 ( .A0(n7627), .A1(n7621), .S(n4049), .Z(n7637) );
  CMX2X1 U16742 ( .A0(n7622), .A1(n7637), .S(n4369), .Z(n7650) );
  CMXI2X1 U16743 ( .A0(n7623), .A1(n7650), .S(n3314), .Z(N2483) );
  CMX2X1 U16744 ( .A0(mem_data1[422]), .A1(mem_data1[423]), .S(n3865), .Z(
        n7633) );
  CMXI2X1 U16745 ( .A0(n7633), .A1(n7624), .S(n4049), .Z(n7640) );
  CMX2X1 U16746 ( .A0(n7625), .A1(n7640), .S(n4369), .Z(n7653) );
  CMXI2X1 U16747 ( .A0(n7626), .A1(n7653), .S(n3482), .Z(N2484) );
  CMX2X1 U16748 ( .A0(mem_data1[423]), .A1(mem_data1[424]), .S(n3877), .Z(
        n7636) );
  CMXI2X1 U16749 ( .A0(n7636), .A1(n7627), .S(n4049), .Z(n7643) );
  CMX2X1 U16750 ( .A0(n7628), .A1(n7643), .S(n4368), .Z(n7656) );
  CMXI2X1 U16751 ( .A0(n7629), .A1(n7656), .S(n3482), .Z(N2485) );
  CMX2X1 U16752 ( .A0(mem_data1[54]), .A1(mem_data1[55]), .S(n3878), .Z(n7696)
         );
  CMXI2X1 U16753 ( .A0(n7696), .A1(n7630), .S(n4049), .Z(n7763) );
  CMX2X1 U16754 ( .A0(n7631), .A1(n7763), .S(n3796), .Z(n7896) );
  CMXI2X1 U16755 ( .A0(n7632), .A1(n7896), .S(n3482), .Z(N2116) );
  CMX2X1 U16756 ( .A0(mem_data1[424]), .A1(mem_data1[425]), .S(n3879), .Z(
        n7639) );
  CMXI2X1 U16757 ( .A0(n7639), .A1(n7633), .S(n4049), .Z(n7646) );
  CMX2X1 U16758 ( .A0(n7634), .A1(n7646), .S(n3776), .Z(n7659) );
  CMXI2X1 U16759 ( .A0(n7635), .A1(n7659), .S(n3482), .Z(N2486) );
  CMX2X1 U16760 ( .A0(mem_data1[425]), .A1(mem_data1[426]), .S(n3880), .Z(
        n7642) );
  CMXI2X1 U16761 ( .A0(n7642), .A1(n7636), .S(n4049), .Z(n7649) );
  CMX2X1 U16762 ( .A0(n7637), .A1(n7649), .S(n4339), .Z(n7662) );
  CMXI2X1 U16763 ( .A0(n7638), .A1(n7662), .S(n3482), .Z(N2487) );
  CMX2X1 U16764 ( .A0(mem_data1[426]), .A1(mem_data1[427]), .S(n3881), .Z(
        n7645) );
  CMXI2X1 U16765 ( .A0(n7645), .A1(n7639), .S(n4049), .Z(n7652) );
  CMX2X1 U16766 ( .A0(n7640), .A1(n7652), .S(n4339), .Z(n7668) );
  CMXI2X1 U16767 ( .A0(n7641), .A1(n7668), .S(n3482), .Z(N2488) );
  CMX2X1 U16768 ( .A0(mem_data1[427]), .A1(mem_data1[428]), .S(n3862), .Z(
        n7648) );
  CMXI2X1 U16769 ( .A0(n7648), .A1(n7642), .S(n4049), .Z(n7655) );
  CMX2X1 U16770 ( .A0(n7643), .A1(n7655), .S(n4339), .Z(n7671) );
  CMXI2X1 U16771 ( .A0(n7644), .A1(n7671), .S(n3482), .Z(N2489) );
  CMX2X1 U16772 ( .A0(mem_data1[428]), .A1(mem_data1[429]), .S(n3863), .Z(
        n7651) );
  CMXI2X1 U16773 ( .A0(n7651), .A1(n7645), .S(n4049), .Z(n7658) );
  CMX2X1 U16774 ( .A0(n7646), .A1(n7658), .S(n4339), .Z(n7674) );
  CMXI2X1 U16775 ( .A0(n7647), .A1(n7674), .S(n3482), .Z(N2490) );
  CMX2X1 U16776 ( .A0(mem_data1[429]), .A1(mem_data1[430]), .S(n3870), .Z(
        n7654) );
  CMXI2X1 U16777 ( .A0(n7654), .A1(n7648), .S(n4049), .Z(n7661) );
  CMX2X1 U16778 ( .A0(n7649), .A1(n7661), .S(n4338), .Z(n7677) );
  CMXI2X1 U16779 ( .A0(n7650), .A1(n7677), .S(n3482), .Z(N2491) );
  CMX2X1 U16780 ( .A0(mem_data1[430]), .A1(mem_data1[431]), .S(n3871), .Z(
        n7657) );
  CMXI2X1 U16781 ( .A0(n7657), .A1(n7651), .S(n4049), .Z(n7667) );
  CMX2X1 U16782 ( .A0(n7652), .A1(n7667), .S(n4338), .Z(n7680) );
  CMXI2X1 U16783 ( .A0(n7653), .A1(n7680), .S(n3481), .Z(N2492) );
  CMX2X1 U16784 ( .A0(mem_data1[431]), .A1(mem_data1[432]), .S(n3864), .Z(
        n7660) );
  CMXI2X1 U16785 ( .A0(n7660), .A1(n7654), .S(n4049), .Z(n7670) );
  CMX2X1 U16786 ( .A0(n7655), .A1(n7670), .S(n4338), .Z(n7683) );
  CMXI2X1 U16787 ( .A0(n7656), .A1(n7683), .S(n3481), .Z(N2493) );
  CMX2X1 U16788 ( .A0(mem_data1[432]), .A1(mem_data1[433]), .S(n3865), .Z(
        n7666) );
  CMXI2X1 U16789 ( .A0(n7666), .A1(n7657), .S(n4049), .Z(n7673) );
  CMX2X1 U16790 ( .A0(n7658), .A1(n7673), .S(n4338), .Z(n7686) );
  CMXI2X1 U16791 ( .A0(n7659), .A1(n7686), .S(n3481), .Z(N2494) );
  CMX2X1 U16792 ( .A0(mem_data1[433]), .A1(mem_data1[434]), .S(n3880), .Z(
        n7669) );
  CMXI2X1 U16793 ( .A0(n7669), .A1(n7660), .S(n4048), .Z(n7676) );
  CMX2X1 U16794 ( .A0(n7661), .A1(n7676), .S(n4338), .Z(n7689) );
  CMXI2X1 U16795 ( .A0(n7662), .A1(n7689), .S(n3481), .Z(N2495) );
  CMX2X1 U16796 ( .A0(mem_data1[55]), .A1(mem_data1[56]), .S(n3881), .Z(n7729)
         );
  CMXI2X1 U16797 ( .A0(n7729), .A1(n7663), .S(n4048), .Z(n7796) );
  CMX2X1 U16798 ( .A0(n7664), .A1(n7796), .S(n4338), .Z(n7929) );
  CMXI2X1 U16799 ( .A0(n7665), .A1(n7929), .S(n3481), .Z(N2117) );
  CMX2X1 U16800 ( .A0(mem_data1[434]), .A1(mem_data1[435]), .S(n3862), .Z(
        n7672) );
  CMXI2X1 U16801 ( .A0(n7672), .A1(n7666), .S(n4048), .Z(n7679) );
  CMX2X1 U16802 ( .A0(n7667), .A1(n7679), .S(n4338), .Z(n7692) );
  CMXI2X1 U16803 ( .A0(n7668), .A1(n7692), .S(n3481), .Z(N2496) );
  CMX2X1 U16804 ( .A0(mem_data1[435]), .A1(mem_data1[436]), .S(n3863), .Z(
        n7675) );
  CMXI2X1 U16805 ( .A0(n7675), .A1(n7669), .S(n4048), .Z(n7682) );
  CMX2X1 U16806 ( .A0(n7670), .A1(n7682), .S(n4338), .Z(n7695) );
  CMXI2X1 U16807 ( .A0(n7671), .A1(n7695), .S(n3481), .Z(N2497) );
  CMX2X1 U16808 ( .A0(mem_data1[436]), .A1(mem_data1[437]), .S(n3873), .Z(
        n7678) );
  CMXI2X1 U16809 ( .A0(n7678), .A1(n7672), .S(n4048), .Z(n7685) );
  CMX2X1 U16810 ( .A0(n7673), .A1(n7685), .S(n4338), .Z(n7701) );
  CMXI2X1 U16811 ( .A0(n7674), .A1(n7701), .S(n3481), .Z(N2498) );
  CMX2X1 U16812 ( .A0(mem_data1[437]), .A1(mem_data1[438]), .S(n3874), .Z(
        n7681) );
  CMXI2X1 U16813 ( .A0(n7681), .A1(n7675), .S(n4048), .Z(n7688) );
  CMX2X1 U16814 ( .A0(n7676), .A1(n7688), .S(n4338), .Z(n7704) );
  CMXI2X1 U16815 ( .A0(n7677), .A1(n7704), .S(n3481), .Z(N2499) );
  CMX2X1 U16816 ( .A0(mem_data1[438]), .A1(mem_data1[439]), .S(n3875), .Z(
        n7684) );
  CMXI2X1 U16817 ( .A0(n7684), .A1(n7678), .S(n4048), .Z(n7691) );
  CMX2X1 U16818 ( .A0(n7679), .A1(n7691), .S(n4338), .Z(n7707) );
  CMXI2X1 U16819 ( .A0(n7680), .A1(n7707), .S(n3484), .Z(N2500) );
  CMX2X1 U16820 ( .A0(mem_data1[439]), .A1(mem_data1[440]), .S(n3876), .Z(
        n7687) );
  CMXI2X1 U16821 ( .A0(n7687), .A1(n7681), .S(n4048), .Z(n7694) );
  CMX2X1 U16822 ( .A0(n7682), .A1(n7694), .S(n4337), .Z(n7710) );
  CMXI2X1 U16823 ( .A0(n7683), .A1(n7710), .S(n3484), .Z(N2501) );
  CMX2X1 U16824 ( .A0(mem_data1[440]), .A1(mem_data1[441]), .S(n3866), .Z(
        n7690) );
  CMXI2X1 U16825 ( .A0(n7690), .A1(n7684), .S(n4048), .Z(n7700) );
  CMX2X1 U16826 ( .A0(n7685), .A1(n7700), .S(n4337), .Z(n7713) );
  CMXI2X1 U16827 ( .A0(n7686), .A1(n7713), .S(n3484), .Z(N2502) );
  CMX2X1 U16828 ( .A0(mem_data1[441]), .A1(mem_data1[442]), .S(n3866), .Z(
        n7693) );
  CMXI2X1 U16829 ( .A0(n7693), .A1(n7687), .S(n4048), .Z(n7703) );
  CMX2X1 U16830 ( .A0(n7688), .A1(n7703), .S(n4337), .Z(n7716) );
  CMXI2X1 U16831 ( .A0(n7689), .A1(n7716), .S(n3526), .Z(N2503) );
  CMX2X1 U16832 ( .A0(mem_data1[442]), .A1(mem_data1[443]), .S(n3867), .Z(
        n7699) );
  CMXI2X1 U16833 ( .A0(n7699), .A1(n7690), .S(n4048), .Z(n7706) );
  CMX2X1 U16834 ( .A0(n7691), .A1(n7706), .S(n4337), .Z(n7719) );
  CMXI2X1 U16835 ( .A0(n7692), .A1(n7719), .S(n3518), .Z(N2504) );
  CMX2X1 U16836 ( .A0(mem_data1[443]), .A1(mem_data1[444]), .S(n3868), .Z(
        n7702) );
  CMXI2X1 U16837 ( .A0(n7702), .A1(n7693), .S(n4048), .Z(n7709) );
  CMX2X1 U16838 ( .A0(n7694), .A1(n7709), .S(n4337), .Z(n7722) );
  CMXI2X1 U16839 ( .A0(n7695), .A1(n7722), .S(n3518), .Z(N2505) );
  CMX2X1 U16840 ( .A0(mem_data1[56]), .A1(mem_data1[57]), .S(n3869), .Z(n7762)
         );
  CMXI2X1 U16841 ( .A0(n7762), .A1(n7696), .S(n4048), .Z(n7829) );
  CMX2X1 U16842 ( .A0(n7697), .A1(n7829), .S(n4337), .Z(n7966) );
  CMXI2X1 U16843 ( .A0(n7698), .A1(n7966), .S(n3518), .Z(N2118) );
  CMX2X1 U16844 ( .A0(mem_data1[444]), .A1(mem_data1[445]), .S(n3870), .Z(
        n7705) );
  CMXI2X1 U16845 ( .A0(n7705), .A1(n7699), .S(n4048), .Z(n7712) );
  CMX2X1 U16846 ( .A0(n7700), .A1(n7712), .S(n4337), .Z(n7725) );
  CMXI2X1 U16847 ( .A0(n7701), .A1(n7725), .S(n3518), .Z(N2506) );
  CMX2X1 U16848 ( .A0(mem_data1[445]), .A1(mem_data1[446]), .S(n3871), .Z(
        n7708) );
  CMXI2X1 U16849 ( .A0(n7708), .A1(n7702), .S(n4048), .Z(n7715) );
  CMX2X1 U16850 ( .A0(n7703), .A1(n7715), .S(n4337), .Z(n7728) );
  CMXI2X1 U16851 ( .A0(n7704), .A1(n7728), .S(n3518), .Z(N2507) );
  CMX2X1 U16852 ( .A0(mem_data1[446]), .A1(mem_data1[447]), .S(n3872), .Z(
        n7711) );
  CMXI2X1 U16853 ( .A0(n7711), .A1(n7705), .S(n4048), .Z(n7718) );
  CMX2X1 U16854 ( .A0(n7706), .A1(n7718), .S(n4337), .Z(n7734) );
  CMXI2X1 U16855 ( .A0(n7707), .A1(n7734), .S(n3518), .Z(N2508) );
  CMX2X1 U16856 ( .A0(mem_data1[447]), .A1(mem_data1[448]), .S(n3872), .Z(
        n7714) );
  CMXI2X1 U16857 ( .A0(n7714), .A1(n7708), .S(n4047), .Z(n7721) );
  CMX2X1 U16858 ( .A0(n7709), .A1(n7721), .S(n4337), .Z(n7737) );
  CMXI2X1 U16859 ( .A0(n7710), .A1(n7737), .S(n3518), .Z(N2509) );
  CMX2X1 U16860 ( .A0(mem_data1[448]), .A1(mem_data1[449]), .S(n3873), .Z(
        n7717) );
  CMXI2X1 U16861 ( .A0(n7717), .A1(n7711), .S(n4047), .Z(n7724) );
  CMX2X1 U16862 ( .A0(n7712), .A1(n7724), .S(n4337), .Z(n7740) );
  CMXI2X1 U16863 ( .A0(n7713), .A1(n7740), .S(n3518), .Z(N2510) );
  CMX2X1 U16864 ( .A0(mem_data1[449]), .A1(mem_data1[450]), .S(n3873), .Z(
        n7720) );
  CMXI2X1 U16865 ( .A0(n7720), .A1(n7714), .S(n4047), .Z(n7727) );
  CMX2X1 U16866 ( .A0(n7715), .A1(n7727), .S(n4336), .Z(n7743) );
  CMXI2X1 U16867 ( .A0(n7716), .A1(n7743), .S(n3517), .Z(N2511) );
  CMX2X1 U16868 ( .A0(mem_data1[450]), .A1(mem_data1[451]), .S(n3874), .Z(
        n7723) );
  CMXI2X1 U16869 ( .A0(n7723), .A1(n7717), .S(n4047), .Z(n7733) );
  CMX2X1 U16870 ( .A0(n7718), .A1(n7733), .S(n4336), .Z(n7746) );
  CMXI2X1 U16871 ( .A0(n7719), .A1(n7746), .S(n3517), .Z(N2512) );
  CMX2X1 U16872 ( .A0(mem_data1[451]), .A1(mem_data1[452]), .S(n3864), .Z(
        n7726) );
  CMXI2X1 U16873 ( .A0(n7726), .A1(n7720), .S(n4047), .Z(n7736) );
  CMX2X1 U16874 ( .A0(n7721), .A1(n7736), .S(n4336), .Z(n7749) );
  CMXI2X1 U16875 ( .A0(n7722), .A1(n7749), .S(n3524), .Z(N2513) );
  CMX2X1 U16876 ( .A0(mem_data1[452]), .A1(mem_data1[453]), .S(n3865), .Z(
        n7732) );
  CMXI2X1 U16877 ( .A0(n7732), .A1(n7723), .S(n4047), .Z(n7739) );
  CMX2X1 U16878 ( .A0(n7724), .A1(n7739), .S(n4336), .Z(n7752) );
  CMXI2X1 U16879 ( .A0(n7725), .A1(n7752), .S(n3517), .Z(N2514) );
  CMX2X1 U16880 ( .A0(mem_data1[453]), .A1(mem_data1[454]), .S(n3866), .Z(
        n7735) );
  CMXI2X1 U16881 ( .A0(n7735), .A1(n7726), .S(n4047), .Z(n7742) );
  CMX2X1 U16882 ( .A0(n7727), .A1(n7742), .S(n4336), .Z(n7755) );
  CMXI2X1 U16883 ( .A0(n7728), .A1(n7755), .S(n3517), .Z(N2515) );
  CMX2X1 U16884 ( .A0(mem_data1[57]), .A1(mem_data1[58]), .S(n3867), .Z(n7795)
         );
  CMXI2X1 U16885 ( .A0(n7795), .A1(n7729), .S(n4047), .Z(n7862) );
  CMX2X1 U16886 ( .A0(n7730), .A1(n7862), .S(n4336), .Z(n7999) );
  CMXI2X1 U16887 ( .A0(n7731), .A1(n7999), .S(n3517), .Z(N2119) );
  CMX2X1 U16888 ( .A0(mem_data1[454]), .A1(mem_data1[455]), .S(n3877), .Z(
        n7738) );
  CMXI2X1 U16889 ( .A0(n7738), .A1(n7732), .S(n4047), .Z(n7745) );
  CMX2X1 U16890 ( .A0(n7733), .A1(n7745), .S(n4336), .Z(n7758) );
  CMXI2X1 U16891 ( .A0(n7734), .A1(n7758), .S(n3517), .Z(N2516) );
  CMX2X1 U16892 ( .A0(mem_data1[455]), .A1(mem_data1[456]), .S(n3878), .Z(
        n7741) );
  CMXI2X1 U16893 ( .A0(n7741), .A1(n7735), .S(n4047), .Z(n7748) );
  CMX2X1 U16894 ( .A0(n7736), .A1(n7748), .S(n4336), .Z(n7761) );
  CMXI2X1 U16895 ( .A0(n7737), .A1(n7761), .S(n3520), .Z(N2517) );
  CMX2X1 U16896 ( .A0(mem_data1[456]), .A1(mem_data1[457]), .S(n3879), .Z(
        n7744) );
  CMXI2X1 U16897 ( .A0(n7744), .A1(n7738), .S(n4047), .Z(n7751) );
  CMX2X1 U16898 ( .A0(n7739), .A1(n7751), .S(n4336), .Z(n7767) );
  CMXI2X1 U16899 ( .A0(n7740), .A1(n7767), .S(n3520), .Z(N2518) );
  CMX2X1 U16900 ( .A0(mem_data1[457]), .A1(mem_data1[458]), .S(n3880), .Z(
        n7747) );
  CMXI2X1 U16901 ( .A0(n7747), .A1(n7741), .S(n4047), .Z(n7754) );
  CMX2X1 U16902 ( .A0(n7742), .A1(n7754), .S(n4336), .Z(n7770) );
  CMXI2X1 U16903 ( .A0(n7743), .A1(n7770), .S(n3520), .Z(N2519) );
  CMX2X1 U16904 ( .A0(mem_data1[458]), .A1(mem_data1[459]), .S(n3867), .Z(
        n7750) );
  CMXI2X1 U16905 ( .A0(n7750), .A1(n7744), .S(n4047), .Z(n7757) );
  CMX2X1 U16906 ( .A0(n7745), .A1(n7757), .S(n4336), .Z(n7773) );
  CMXI2X1 U16907 ( .A0(n7746), .A1(n7773), .S(n3520), .Z(N2520) );
  CMX2X1 U16908 ( .A0(mem_data1[459]), .A1(mem_data1[460]), .S(n3875), .Z(
        n7753) );
  CMXI2X1 U16909 ( .A0(n7753), .A1(n7747), .S(n4047), .Z(n7760) );
  CMX2X1 U16910 ( .A0(n7748), .A1(n7760), .S(n4335), .Z(n7776) );
  CMXI2X1 U16911 ( .A0(n7749), .A1(n7776), .S(n3520), .Z(N2521) );
  CMX2X1 U16912 ( .A0(mem_data1[460]), .A1(mem_data1[461]), .S(n3876), .Z(
        n7756) );
  CMXI2X1 U16913 ( .A0(n7756), .A1(n7750), .S(n4047), .Z(n7766) );
  CMX2X1 U16914 ( .A0(n7751), .A1(n7766), .S(n4335), .Z(n7779) );
  CMXI2X1 U16915 ( .A0(n7752), .A1(n7779), .S(n3520), .Z(N2522) );
  CMX2X1 U16916 ( .A0(mem_data1[461]), .A1(mem_data1[462]), .S(n3877), .Z(
        n7759) );
  CMXI2X1 U16917 ( .A0(n7759), .A1(n7753), .S(n4047), .Z(n7769) );
  CMX2X1 U16918 ( .A0(n7754), .A1(n7769), .S(n4335), .Z(n7782) );
  CMXI2X1 U16919 ( .A0(n7755), .A1(n7782), .S(n3520), .Z(N2523) );
  CMX2X1 U16920 ( .A0(mem_data1[462]), .A1(mem_data1[463]), .S(n3878), .Z(
        n7765) );
  CMXI2X1 U16921 ( .A0(n7765), .A1(n7756), .S(n4046), .Z(n7772) );
  CMX2X1 U16922 ( .A0(n7757), .A1(n7772), .S(n4335), .Z(n7785) );
  CMXI2X1 U16923 ( .A0(n7758), .A1(n7785), .S(n3519), .Z(N2524) );
  CMX2X1 U16924 ( .A0(mem_data1[463]), .A1(mem_data1[464]), .S(n3879), .Z(
        n7768) );
  CMXI2X1 U16925 ( .A0(n7768), .A1(n7759), .S(n4046), .Z(n7775) );
  CMX2X1 U16926 ( .A0(n7760), .A1(n7775), .S(n4335), .Z(n7788) );
  CMXI2X1 U16927 ( .A0(n7761), .A1(n7788), .S(n3519), .Z(N2525) );
  CMX2X1 U16928 ( .A0(mem_data1[58]), .A1(mem_data1[59]), .S(n3880), .Z(n7828)
         );
  CMXI2X1 U16929 ( .A0(n7828), .A1(n7762), .S(n4046), .Z(n7895) );
  CMX2X1 U16930 ( .A0(n7763), .A1(n7895), .S(n4335), .Z(n8032) );
  CMXI2X1 U16931 ( .A0(n7764), .A1(n8032), .S(n3519), .Z(N2120) );
  CMX2X1 U16932 ( .A0(mem_data1[464]), .A1(mem_data1[465]), .S(n3881), .Z(
        n7771) );
  CMXI2X1 U16933 ( .A0(n7771), .A1(n7765), .S(n4046), .Z(n7778) );
  CMX2X1 U16934 ( .A0(n7766), .A1(n7778), .S(n4335), .Z(n7791) );
  CMXI2X1 U16935 ( .A0(n7767), .A1(n7791), .S(n3519), .Z(N2526) );
  CMX2X1 U16936 ( .A0(mem_data1[465]), .A1(mem_data1[466]), .S(n3874), .Z(
        n7774) );
  CMXI2X1 U16937 ( .A0(n7774), .A1(n7768), .S(n4046), .Z(n7781) );
  CMX2X1 U16938 ( .A0(n7769), .A1(n7781), .S(n4335), .Z(n7794) );
  CMXI2X1 U16939 ( .A0(n7770), .A1(n7794), .S(n3519), .Z(N2527) );
  CMX2X1 U16940 ( .A0(mem_data1[466]), .A1(mem_data1[467]), .S(n3875), .Z(
        n7777) );
  CMXI2X1 U16941 ( .A0(n7777), .A1(n7771), .S(n4046), .Z(n7784) );
  CMX2X1 U16942 ( .A0(n7772), .A1(n7784), .S(n4335), .Z(n7800) );
  CMXI2X1 U16943 ( .A0(n7773), .A1(n7800), .S(n3519), .Z(N2528) );
  CMX2X1 U16944 ( .A0(mem_data1[467]), .A1(mem_data1[468]), .S(n3862), .Z(
        n7780) );
  CMXI2X1 U16945 ( .A0(n7780), .A1(n7774), .S(n4046), .Z(n7787) );
  CMX2X1 U16946 ( .A0(n7775), .A1(n7787), .S(n4335), .Z(n7803) );
  CMXI2X1 U16947 ( .A0(n7776), .A1(n7803), .S(n3519), .Z(N2529) );
  CMX2X1 U16948 ( .A0(mem_data1[468]), .A1(mem_data1[469]), .S(n3863), .Z(
        n7783) );
  CMXI2X1 U16949 ( .A0(n7783), .A1(n7777), .S(n4046), .Z(n7790) );
  CMX2X1 U16950 ( .A0(n7778), .A1(n7790), .S(n4335), .Z(n7806) );
  CMXI2X1 U16951 ( .A0(n7779), .A1(n7806), .S(n3519), .Z(N2530) );
  CMX2X1 U16952 ( .A0(mem_data1[469]), .A1(mem_data1[470]), .S(n3868), .Z(
        n7786) );
  CMXI2X1 U16953 ( .A0(n7786), .A1(n7780), .S(n4046), .Z(n7793) );
  CMX2X1 U16954 ( .A0(n7781), .A1(n7793), .S(n4334), .Z(n7809) );
  CMXI2X1 U16955 ( .A0(n7782), .A1(n7809), .S(n3519), .Z(N2531) );
  CMX2X1 U16956 ( .A0(mem_data1[470]), .A1(mem_data1[471]), .S(n3869), .Z(
        n7789) );
  CMXI2X1 U16957 ( .A0(n7789), .A1(n7783), .S(n4046), .Z(n7799) );
  CMX2X1 U16958 ( .A0(n7784), .A1(n7799), .S(n4334), .Z(n7812) );
  CMXI2X1 U16959 ( .A0(n7785), .A1(n7812), .S(n3519), .Z(N2532) );
  CMX2X1 U16960 ( .A0(mem_data1[471]), .A1(mem_data1[472]), .S(n3870), .Z(
        n7792) );
  CMXI2X1 U16961 ( .A0(n7792), .A1(n7786), .S(n4046), .Z(n7802) );
  CMX2X1 U16962 ( .A0(n7787), .A1(n7802), .S(n4334), .Z(n7815) );
  CMXI2X1 U16963 ( .A0(n7788), .A1(n7815), .S(n3519), .Z(N2533) );
  CMX2X1 U16964 ( .A0(mem_data1[472]), .A1(mem_data1[473]), .S(n3871), .Z(
        n7798) );
  CMXI2X1 U16965 ( .A0(n7798), .A1(n7789), .S(n4046), .Z(n7805) );
  CMX2X1 U16966 ( .A0(n7790), .A1(n7805), .S(n4334), .Z(n7818) );
  CMXI2X1 U16967 ( .A0(n7791), .A1(n7818), .S(n3522), .Z(N2534) );
  CMX2X1 U16968 ( .A0(mem_data1[473]), .A1(mem_data1[474]), .S(n3881), .Z(
        n7801) );
  CMXI2X1 U16969 ( .A0(n7801), .A1(n7792), .S(n4046), .Z(n7808) );
  CMX2X1 U16970 ( .A0(n7793), .A1(n7808), .S(n4334), .Z(n7821) );
  CMXI2X1 U16971 ( .A0(n7794), .A1(n7821), .S(n3522), .Z(N2535) );
  CMX2X1 U16972 ( .A0(mem_data1[59]), .A1(mem_data1[60]), .S(n3862), .Z(n7861)
         );
  CMXI2X1 U16973 ( .A0(n7861), .A1(n7795), .S(n4046), .Z(n7928) );
  CMX2X1 U16974 ( .A0(n7796), .A1(n7928), .S(n4334), .Z(n8065) );
  CMXI2X1 U16975 ( .A0(n7797), .A1(n8065), .S(n3522), .Z(N2121) );
  CMX2X1 U16976 ( .A0(mem_data1[474]), .A1(mem_data1[475]), .S(n3863), .Z(
        n7804) );
  CMXI2X1 U16977 ( .A0(n7804), .A1(n7798), .S(n4046), .Z(n7811) );
  CMX2X1 U16978 ( .A0(n7799), .A1(n7811), .S(n4334), .Z(n7824) );
  CMXI2X1 U16979 ( .A0(n7800), .A1(n7824), .S(n3521), .Z(N2536) );
  CMX2X1 U16980 ( .A0(mem_data1[475]), .A1(mem_data1[476]), .S(n3864), .Z(
        n7807) );
  CMXI2X1 U16981 ( .A0(n7807), .A1(n7801), .S(n4046), .Z(n7814) );
  CMX2X1 U16982 ( .A0(n7802), .A1(n7814), .S(n4334), .Z(n7827) );
  CMXI2X1 U16983 ( .A0(n7803), .A1(n7827), .S(n3521), .Z(N2537) );
  CMX2X1 U16984 ( .A0(mem_data1[476]), .A1(mem_data1[477]), .S(n3868), .Z(
        n7810) );
  CMXI2X1 U16985 ( .A0(n7810), .A1(n7804), .S(n4045), .Z(n7817) );
  CMX2X1 U16986 ( .A0(n7805), .A1(n7817), .S(n4334), .Z(n7833) );
  CMXI2X1 U16987 ( .A0(n7806), .A1(n7833), .S(n3521), .Z(N2538) );
  CMX2X1 U16988 ( .A0(mem_data1[477]), .A1(mem_data1[478]), .S(n3864), .Z(
        n7813) );
  CMXI2X1 U16989 ( .A0(n7813), .A1(n7807), .S(n4045), .Z(n7820) );
  CMX2X1 U16990 ( .A0(n7808), .A1(n7820), .S(n4334), .Z(n7836) );
  CMXI2X1 U16991 ( .A0(n7809), .A1(n7836), .S(n3521), .Z(N2539) );
  CMX2X1 U16992 ( .A0(mem_data1[478]), .A1(mem_data1[479]), .S(n3865), .Z(
        n7816) );
  CMXI2X1 U16993 ( .A0(n7816), .A1(n7810), .S(n4045), .Z(n7823) );
  CMX2X1 U16994 ( .A0(n7811), .A1(n7823), .S(n4334), .Z(n7839) );
  CMXI2X1 U16995 ( .A0(n7812), .A1(n7839), .S(n3521), .Z(N2540) );
  CMX2X1 U16996 ( .A0(mem_data1[479]), .A1(mem_data1[480]), .S(n3866), .Z(
        n7819) );
  CMXI2X1 U16997 ( .A0(n7819), .A1(n7813), .S(n4045), .Z(n7826) );
  CMX2X1 U16998 ( .A0(n7814), .A1(n7826), .S(n4333), .Z(n7842) );
  CMXI2X1 U16999 ( .A0(n7815), .A1(n7842), .S(n3521), .Z(N2541) );
  CMX2X1 U17000 ( .A0(mem_data1[480]), .A1(mem_data1[481]), .S(n3867), .Z(
        n7822) );
  CMXI2X1 U17001 ( .A0(n7822), .A1(n7816), .S(n4045), .Z(n7832) );
  CMX2X1 U17002 ( .A0(n7817), .A1(n7832), .S(n4333), .Z(n7845) );
  CMXI2X1 U17003 ( .A0(n7818), .A1(n7845), .S(n3521), .Z(N2542) );
  CMX2X1 U17004 ( .A0(mem_data1[481]), .A1(mem_data1[482]), .S(n3868), .Z(
        n7825) );
  CMXI2X1 U17005 ( .A0(n7825), .A1(n7819), .S(n4045), .Z(n7835) );
  CMX2X1 U17006 ( .A0(n7820), .A1(n7835), .S(n4333), .Z(n7848) );
  CMXI2X1 U17007 ( .A0(n7821), .A1(n7848), .S(n3521), .Z(N2543) );
  CMX2X1 U17008 ( .A0(mem_data1[482]), .A1(mem_data1[483]), .S(n3869), .Z(
        n7831) );
  CMXI2X1 U17009 ( .A0(n7831), .A1(n7822), .S(n4045), .Z(n7838) );
  CMX2X1 U17010 ( .A0(n7823), .A1(n7838), .S(n4333), .Z(n7851) );
  CMXI2X1 U17011 ( .A0(n7824), .A1(n7851), .S(n3521), .Z(N2544) );
  CMX2X1 U17012 ( .A0(mem_data1[483]), .A1(mem_data1[484]), .S(n3870), .Z(
        n7834) );
  CMXI2X1 U17013 ( .A0(n7834), .A1(n7825), .S(n4045), .Z(n7841) );
  CMX2X1 U17014 ( .A0(n7826), .A1(n7841), .S(n4333), .Z(n7854) );
  CMXI2X1 U17015 ( .A0(n7827), .A1(n7854), .S(n3521), .Z(N2545) );
  CMX2X1 U17016 ( .A0(mem_data1[60]), .A1(mem_data1[61]), .S(n3876), .Z(n7894)
         );
  CMXI2X1 U17017 ( .A0(n7894), .A1(n7828), .S(n4045), .Z(n7965) );
  CMX2X1 U17018 ( .A0(n7829), .A1(n7965), .S(n4333), .Z(n8098) );
  CMXI2X1 U17019 ( .A0(n7830), .A1(n8098), .S(n3521), .Z(N2122) );
  CMX2X1 U17020 ( .A0(mem_data1[484]), .A1(mem_data1[485]), .S(n3877), .Z(
        n7837) );
  CMXI2X1 U17021 ( .A0(n7837), .A1(n7831), .S(n4045), .Z(n7844) );
  CMX2X1 U17022 ( .A0(n7832), .A1(n7844), .S(n4333), .Z(n7857) );
  CMXI2X1 U17023 ( .A0(n7833), .A1(n7857), .S(n3520), .Z(N2546) );
  CMX2X1 U17024 ( .A0(mem_data1[485]), .A1(mem_data1[486]), .S(n3871), .Z(
        n7840) );
  CMXI2X1 U17025 ( .A0(n7840), .A1(n7834), .S(n4045), .Z(n7847) );
  CMX2X1 U17026 ( .A0(n7835), .A1(n7847), .S(n4333), .Z(n7860) );
  CMXI2X1 U17027 ( .A0(n7836), .A1(n7860), .S(n3520), .Z(N2547) );
  CMX2X1 U17028 ( .A0(mem_data1[486]), .A1(mem_data1[487]), .S(n3872), .Z(
        n7843) );
  CMXI2X1 U17029 ( .A0(n7843), .A1(n7837), .S(n4045), .Z(n7850) );
  CMX2X1 U17030 ( .A0(n7838), .A1(n7850), .S(n4333), .Z(n7866) );
  CMXI2X1 U17031 ( .A0(n7839), .A1(n7866), .S(n3520), .Z(N2548) );
  CMX2X1 U17032 ( .A0(mem_data1[487]), .A1(mem_data1[488]), .S(n3872), .Z(
        n7846) );
  CMXI2X1 U17033 ( .A0(n7846), .A1(n7840), .S(n4045), .Z(n7853) );
  CMX2X1 U17034 ( .A0(n7841), .A1(n7853), .S(n4333), .Z(n7869) );
  CMXI2X1 U17035 ( .A0(n7842), .A1(n7869), .S(n3520), .Z(N2549) );
  CMX2X1 U17036 ( .A0(mem_data1[488]), .A1(mem_data1[489]), .S(n3873), .Z(
        n7849) );
  CMXI2X1 U17037 ( .A0(n7849), .A1(n7843), .S(n4045), .Z(n7856) );
  CMX2X1 U17038 ( .A0(n7844), .A1(n7856), .S(n4333), .Z(n7872) );
  CMXI2X1 U17039 ( .A0(n7845), .A1(n7872), .S(n3523), .Z(N2550) );
  CMX2X1 U17040 ( .A0(mem_data1[489]), .A1(mem_data1[490]), .S(n3874), .Z(
        n7852) );
  CMXI2X1 U17041 ( .A0(n7852), .A1(n7846), .S(n4045), .Z(n7859) );
  CMX2X1 U17042 ( .A0(n7847), .A1(n7859), .S(n4332), .Z(n7875) );
  CMXI2X1 U17043 ( .A0(n7848), .A1(n7875), .S(n3523), .Z(N2551) );
  CMX2X1 U17044 ( .A0(mem_data1[490]), .A1(mem_data1[491]), .S(n3875), .Z(
        n7855) );
  CMXI2X1 U17045 ( .A0(n7855), .A1(n7849), .S(n4045), .Z(n7865) );
  CMX2X1 U17046 ( .A0(n7850), .A1(n7865), .S(n4332), .Z(n7878) );
  CMXI2X1 U17047 ( .A0(n7851), .A1(n7878), .S(n3523), .Z(N2552) );
  CMX2X1 U17048 ( .A0(mem_data1[491]), .A1(mem_data1[492]), .S(n3865), .Z(
        n7858) );
  CMXI2X1 U17049 ( .A0(n7858), .A1(n7852), .S(n4044), .Z(n7868) );
  CMX2X1 U17050 ( .A0(n7853), .A1(n7868), .S(n4332), .Z(n7881) );
  CMXI2X1 U17051 ( .A0(n7854), .A1(n7881), .S(n3523), .Z(N2553) );
  CMX2X1 U17052 ( .A0(mem_data1[492]), .A1(mem_data1[493]), .S(n3866), .Z(
        n7864) );
  CMXI2X1 U17053 ( .A0(n7864), .A1(n7855), .S(n4044), .Z(n7871) );
  CMX2X1 U17054 ( .A0(n7856), .A1(n7871), .S(n4332), .Z(n7884) );
  CMXI2X1 U17055 ( .A0(n7857), .A1(n7884), .S(n3523), .Z(N2554) );
  CMX2X1 U17056 ( .A0(mem_data1[493]), .A1(mem_data1[494]), .S(n3867), .Z(
        n7867) );
  CMXI2X1 U17057 ( .A0(n7867), .A1(n7858), .S(n4044), .Z(n7874) );
  CMX2X1 U17058 ( .A0(n7859), .A1(n7874), .S(n4332), .Z(n7887) );
  CMXI2X1 U17059 ( .A0(n7860), .A1(n7887), .S(n3523), .Z(N2555) );
  CMX2X1 U17060 ( .A0(mem_data1[61]), .A1(mem_data1[62]), .S(n3868), .Z(n7927)
         );
  CMXI2X1 U17061 ( .A0(n7927), .A1(n7861), .S(n4044), .Z(n7998) );
  CMX2X1 U17062 ( .A0(n7862), .A1(n7998), .S(n4332), .Z(n8131) );
  CMXI2X1 U17063 ( .A0(n7863), .A1(n8131), .S(n3523), .Z(N2123) );
  CMX2X1 U17064 ( .A0(mem_data1[494]), .A1(mem_data1[495]), .S(n3869), .Z(
        n7870) );
  CMXI2X1 U17065 ( .A0(n7870), .A1(n7864), .S(n4044), .Z(n7877) );
  CMX2X1 U17066 ( .A0(n7865), .A1(n7877), .S(n4332), .Z(n7890) );
  CMXI2X1 U17067 ( .A0(n7866), .A1(n7890), .S(n3523), .Z(N2556) );
  CMX2X1 U17068 ( .A0(mem_data1[495]), .A1(mem_data1[496]), .S(n3873), .Z(
        n7873) );
  CMXI2X1 U17069 ( .A0(n7873), .A1(n7867), .S(n4044), .Z(n7880) );
  CMX2X1 U17070 ( .A0(n7868), .A1(n7880), .S(n4332), .Z(n7893) );
  CMXI2X1 U17071 ( .A0(n7869), .A1(n7893), .S(n3523), .Z(N2557) );
  CMX2X1 U17072 ( .A0(mem_data1[496]), .A1(mem_data1[497]), .S(n3874), .Z(
        n7876) );
  CMXI2X1 U17073 ( .A0(n7876), .A1(n7870), .S(n4044), .Z(n7883) );
  CMX2X1 U17074 ( .A0(n7871), .A1(n7883), .S(n4332), .Z(n7899) );
  CMXI2X1 U17075 ( .A0(n7872), .A1(n7899), .S(n3523), .Z(N2558) );
  CMX2X1 U17076 ( .A0(mem_data1[497]), .A1(mem_data1[498]), .S(n3875), .Z(
        n7879) );
  CMXI2X1 U17077 ( .A0(n7879), .A1(n7873), .S(n4044), .Z(n7886) );
  CMX2X1 U17078 ( .A0(n7874), .A1(n7886), .S(n4332), .Z(n7902) );
  CMXI2X1 U17079 ( .A0(n7875), .A1(n7902), .S(n3522), .Z(N2559) );
  CMX2X1 U17080 ( .A0(mem_data1[498]), .A1(mem_data1[499]), .S(n3876), .Z(
        n7882) );
  CMXI2X1 U17081 ( .A0(n7882), .A1(n7876), .S(n4044), .Z(n7889) );
  CMX2X1 U17082 ( .A0(n7877), .A1(n7889), .S(n4332), .Z(n7905) );
  CMXI2X1 U17083 ( .A0(n7878), .A1(n7905), .S(n3522), .Z(N2560) );
  CMX2X1 U17084 ( .A0(mem_data1[499]), .A1(mem_data1[500]), .S(n3877), .Z(
        n7885) );
  CMXI2X1 U17085 ( .A0(n7885), .A1(n7879), .S(n4044), .Z(n7892) );
  CMX2X1 U17086 ( .A0(n7880), .A1(n7892), .S(n4331), .Z(n7908) );
  CMXI2X1 U17087 ( .A0(n7881), .A1(n7908), .S(n3522), .Z(N2561) );
  CMX2X1 U17088 ( .A0(mem_data1[500]), .A1(mem_data1[501]), .S(n3879), .Z(
        n7888) );
  CMXI2X1 U17089 ( .A0(n7888), .A1(n7882), .S(n4044), .Z(n7898) );
  CMX2X1 U17090 ( .A0(n7883), .A1(n7898), .S(n4331), .Z(n7911) );
  CMXI2X1 U17091 ( .A0(n7884), .A1(n7911), .S(n3522), .Z(N2562) );
  CMX2X1 U17092 ( .A0(mem_data1[501]), .A1(mem_data1[502]), .S(n3878), .Z(
        n7891) );
  CMXI2X1 U17093 ( .A0(n7891), .A1(n7885), .S(n4044), .Z(n7901) );
  CMX2X1 U17094 ( .A0(n7886), .A1(n7901), .S(n4331), .Z(n7914) );
  CMXI2X1 U17095 ( .A0(n7887), .A1(n7914), .S(n3522), .Z(N2563) );
  CMX2X1 U17096 ( .A0(mem_data1[502]), .A1(mem_data1[503]), .S(n3879), .Z(
        n7897) );
  CMXI2X1 U17097 ( .A0(n7897), .A1(n7888), .S(n4044), .Z(n7904) );
  CMX2X1 U17098 ( .A0(n7889), .A1(n7904), .S(n4331), .Z(n7917) );
  CMXI2X1 U17099 ( .A0(n7890), .A1(n7917), .S(n3522), .Z(N2564) );
  CMX2X1 U17100 ( .A0(mem_data1[503]), .A1(mem_data1[504]), .S(n3880), .Z(
        n7900) );
  CMXI2X1 U17101 ( .A0(n7900), .A1(n7891), .S(n4044), .Z(n7907) );
  CMX2X1 U17102 ( .A0(n7892), .A1(n7907), .S(n4331), .Z(n7920) );
  CMXI2X1 U17103 ( .A0(n7893), .A1(n7920), .S(n3522), .Z(N2565) );
  CMX2X1 U17104 ( .A0(mem_data1[62]), .A1(mem_data1[63]), .S(n3866), .Z(n7964)
         );
  CMXI2X1 U17105 ( .A0(n7964), .A1(n7894), .S(n4044), .Z(n8031) );
  CMX2X1 U17106 ( .A0(n7895), .A1(n8031), .S(n4331), .Z(n8164) );
  CMXI2X1 U17107 ( .A0(n7896), .A1(n8164), .S(n3522), .Z(N2124) );
  CMX2X1 U17108 ( .A0(mem_data1[504]), .A1(mem_data1[505]), .S(n3867), .Z(
        n7903) );
  CMXI2X1 U17109 ( .A0(n7903), .A1(n7897), .S(n4044), .Z(n7910) );
  CMX2X1 U17110 ( .A0(n7898), .A1(n7910), .S(n4331), .Z(n7923) );
  CMXI2X1 U17111 ( .A0(n7899), .A1(n7923), .S(n3525), .Z(N2566) );
  CMX2X1 U17112 ( .A0(mem_data1[505]), .A1(mem_data1[506]), .S(n3868), .Z(
        n7906) );
  CMXI2X1 U17113 ( .A0(n7906), .A1(n7900), .S(n4043), .Z(n7913) );
  CMX2X1 U17114 ( .A0(n7901), .A1(n7913), .S(n4331), .Z(n7926) );
  CMXI2X1 U17115 ( .A0(n7902), .A1(n7926), .S(n3525), .Z(N2567) );
  CMX2X1 U17116 ( .A0(mem_data1[506]), .A1(mem_data1[507]), .S(n3864), .Z(
        n7909) );
  CMXI2X1 U17117 ( .A0(n7909), .A1(n7903), .S(n4043), .Z(n7916) );
  CMX2X1 U17118 ( .A0(n7904), .A1(n7916), .S(n4331), .Z(n7936) );
  CMXI2X1 U17119 ( .A0(n7905), .A1(n7936), .S(n3525), .Z(N2568) );
  CMX2X1 U17120 ( .A0(mem_data1[507]), .A1(mem_data1[508]), .S(n3865), .Z(
        n7912) );
  CMXI2X1 U17121 ( .A0(n7912), .A1(n7906), .S(n4043), .Z(n7919) );
  CMX2X1 U17122 ( .A0(n7907), .A1(n7919), .S(n4331), .Z(n7939) );
  CMXI2X1 U17123 ( .A0(n7908), .A1(n7939), .S(n3525), .Z(N2569) );
  CMX2X1 U17124 ( .A0(mem_data1[508]), .A1(mem_data1[509]), .S(n3869), .Z(
        n7915) );
  CMXI2X1 U17125 ( .A0(n7915), .A1(n7909), .S(n4043), .Z(n7922) );
  CMX2X1 U17126 ( .A0(n7910), .A1(n7922), .S(n4331), .Z(n7942) );
  CMXI2X1 U17127 ( .A0(n7911), .A1(n7942), .S(n3525), .Z(N2570) );
  CMX2X1 U17128 ( .A0(mem_data1[509]), .A1(mem_data1[510]), .S(n3870), .Z(
        n7918) );
  CMXI2X1 U17129 ( .A0(n7918), .A1(n7912), .S(n4043), .Z(n7925) );
  CMX2X1 U17130 ( .A0(n7913), .A1(n7925), .S(n4330), .Z(n7945) );
  CMXI2X1 U17131 ( .A0(n7914), .A1(n7945), .S(n3525), .Z(N2571) );
  CMX2X1 U17132 ( .A0(mem_data1[510]), .A1(mem_data1[511]), .S(n3872), .Z(
        n7921) );
  CMXI2X1 U17133 ( .A0(n7921), .A1(n7915), .S(n4043), .Z(n7935) );
  CMX2X1 U17134 ( .A0(n7916), .A1(n7935), .S(n4330), .Z(n7948) );
  CMXI2X1 U17135 ( .A0(n7917), .A1(n7948), .S(n3525), .Z(N2572) );
  CMX2X1 U17136 ( .A0(mem_data1[511]), .A1(mem_data1[512]), .S(n3873), .Z(
        n7924) );
  CMXI2X1 U17137 ( .A0(n7924), .A1(n7918), .S(n4043), .Z(n7938) );
  CMX2X1 U17138 ( .A0(n7919), .A1(n7938), .S(n4330), .Z(n7951) );
  CMXI2X1 U17139 ( .A0(n7920), .A1(n7951), .S(n3524), .Z(N2573) );
  CMX2X1 U17140 ( .A0(mem_data1[512]), .A1(mem_data1[513]), .S(n3874), .Z(
        n7934) );
  CMXI2X1 U17141 ( .A0(n7934), .A1(n7921), .S(n4043), .Z(n7941) );
  CMX2X1 U17142 ( .A0(n7922), .A1(n7941), .S(n4330), .Z(n7954) );
  CMXI2X1 U17143 ( .A0(n7923), .A1(n7954), .S(n3524), .Z(N2574) );
  CMX2X1 U17144 ( .A0(mem_data1[513]), .A1(mem_data1[514]), .S(n3875), .Z(
        n7937) );
  CMXI2X1 U17145 ( .A0(n7937), .A1(n7924), .S(n4043), .Z(n7944) );
  CMX2X1 U17146 ( .A0(n7925), .A1(n7944), .S(n4330), .Z(n7957) );
  CMXI2X1 U17147 ( .A0(n7926), .A1(n7957), .S(n3524), .Z(N2575) );
  CMX2X1 U17148 ( .A0(mem_data1[63]), .A1(mem_data1[64]), .S(n3872), .Z(n7997)
         );
  CMXI2X1 U17149 ( .A0(n7997), .A1(n7927), .S(n4043), .Z(n8064) );
  CMX2X1 U17150 ( .A0(n7928), .A1(n8064), .S(n4330), .Z(n8197) );
  CMXI2X1 U17151 ( .A0(n7929), .A1(n8197), .S(n3524), .Z(N2125) );
  CMXI2X1 U17152 ( .A0(n4416), .A1(n7931), .S(n3783), .Z(n7933) );
  CMXI2X1 U17153 ( .A0(n7933), .A1(n7932), .S(n3524), .Z(N2080) );
  CMX2X1 U17154 ( .A0(mem_data1[514]), .A1(mem_data1[515]), .S(n3873), .Z(
        n7940) );
  CMXI2X1 U17155 ( .A0(n7940), .A1(n7934), .S(n4043), .Z(n7947) );
  CMX2X1 U17156 ( .A0(n7935), .A1(n7947), .S(n4330), .Z(n7960) );
  CMXI2X1 U17157 ( .A0(n7936), .A1(n7960), .S(n3524), .Z(N2576) );
  CMX2X1 U17158 ( .A0(mem_data1[515]), .A1(mem_data1[516]), .S(n3874), .Z(
        n7943) );
  CMXI2X1 U17159 ( .A0(n7943), .A1(n7937), .S(n4043), .Z(n7950) );
  CMX2X1 U17160 ( .A0(n7938), .A1(n7950), .S(n4330), .Z(n7963) );
  CMXI2X1 U17161 ( .A0(n7939), .A1(n7963), .S(n3524), .Z(N2577) );
  CMX2X1 U17162 ( .A0(mem_data1[516]), .A1(mem_data1[517]), .S(n3875), .Z(
        n7946) );
  CMXI2X1 U17163 ( .A0(n7946), .A1(n7940), .S(n4043), .Z(n7953) );
  CMX2X1 U17164 ( .A0(n7941), .A1(n7953), .S(n4330), .Z(n7969) );
  CMXI2X1 U17165 ( .A0(n7942), .A1(n7969), .S(n3524), .Z(N2578) );
  CMX2X1 U17166 ( .A0(mem_data1[517]), .A1(mem_data1[518]), .S(n3874), .Z(
        n7949) );
  CMXI2X1 U17167 ( .A0(n7949), .A1(n7943), .S(n4043), .Z(n7956) );
  CMX2X1 U17168 ( .A0(n7944), .A1(n7956), .S(n4330), .Z(n7972) );
  CMXI2X1 U17169 ( .A0(n7945), .A1(n7972), .S(n3524), .Z(N2579) );
  CMX2X1 U17170 ( .A0(mem_data1[518]), .A1(mem_data1[519]), .S(n3871), .Z(
        n7952) );
  CMXI2X1 U17171 ( .A0(n7952), .A1(n7946), .S(n4043), .Z(n7959) );
  CMX2X1 U17172 ( .A0(n7947), .A1(n7959), .S(n4329), .Z(n7975) );
  CMXI2X1 U17173 ( .A0(n7948), .A1(n7975), .S(n3524), .Z(N2580) );
  CMX2X1 U17174 ( .A0(mem_data1[519]), .A1(mem_data1[520]), .S(n3872), .Z(
        n7955) );
  CMXI2X1 U17175 ( .A0(n7955), .A1(n7949), .S(n4043), .Z(n7962) );
  CMX2X1 U17176 ( .A0(n7950), .A1(n7962), .S(n4329), .Z(n7978) );
  CMXI2X1 U17177 ( .A0(n7951), .A1(n7978), .S(n3523), .Z(N2581) );
  CMX2X1 U17178 ( .A0(mem_data1[520]), .A1(mem_data1[521]), .S(n3873), .Z(
        n7958) );
  CMXI2X1 U17179 ( .A0(n7958), .A1(n7952), .S(n4042), .Z(n7968) );
  CMX2X1 U17180 ( .A0(n7953), .A1(n7968), .S(n4329), .Z(n7981) );
  CMXI2X1 U17181 ( .A0(n7954), .A1(n7981), .S(n3527), .Z(N2582) );
  CMX2X1 U17182 ( .A0(mem_data1[521]), .A1(mem_data1[522]), .S(n3874), .Z(
        n7961) );
  CMXI2X1 U17183 ( .A0(n7961), .A1(n7955), .S(n4042), .Z(n7971) );
  CMX2X1 U17184 ( .A0(n7956), .A1(n7971), .S(n4329), .Z(n7984) );
  CMXI2X1 U17185 ( .A0(n7957), .A1(n7984), .S(n3527), .Z(N2583) );
  CMX2X1 U17186 ( .A0(mem_data1[522]), .A1(mem_data1[523]), .S(n3875), .Z(
        n7967) );
  CMXI2X1 U17187 ( .A0(n7967), .A1(n7958), .S(n4042), .Z(n7974) );
  CMX2X1 U17188 ( .A0(n7959), .A1(n7974), .S(n4329), .Z(n7987) );
  CMXI2X1 U17189 ( .A0(n7960), .A1(n7987), .S(n3527), .Z(N2584) );
  CMX2X1 U17190 ( .A0(mem_data1[523]), .A1(mem_data1[524]), .S(n3876), .Z(
        n7970) );
  CMXI2X1 U17191 ( .A0(n7970), .A1(n7961), .S(n4042), .Z(n7977) );
  CMX2X1 U17192 ( .A0(n7962), .A1(n7977), .S(n4329), .Z(n7990) );
  CMXI2X1 U17193 ( .A0(n7963), .A1(n7990), .S(n3526), .Z(N2585) );
  CMX2X1 U17194 ( .A0(mem_data1[64]), .A1(mem_data1[65]), .S(n3881), .Z(n8030)
         );
  CMXI2X1 U17195 ( .A0(n8030), .A1(n7964), .S(n4042), .Z(n8097) );
  CMX2X1 U17196 ( .A0(n7965), .A1(n8097), .S(n4329), .Z(n8230) );
  CMXI2X1 U17197 ( .A0(n7966), .A1(n8230), .S(n3526), .Z(N2126) );
  CMX2X1 U17198 ( .A0(mem_data1[524]), .A1(mem_data1[525]), .S(n3876), .Z(
        n7973) );
  CMXI2X1 U17199 ( .A0(n7973), .A1(n7967), .S(n4042), .Z(n7980) );
  CMX2X1 U17200 ( .A0(n7968), .A1(n7980), .S(n4329), .Z(n7993) );
  CMXI2X1 U17201 ( .A0(n7969), .A1(n7993), .S(n3526), .Z(N2586) );
  CMX2X1 U17202 ( .A0(mem_data1[525]), .A1(mem_data1[526]), .S(n3877), .Z(
        n7976) );
  CMXI2X1 U17203 ( .A0(n7976), .A1(n7970), .S(n4042), .Z(n7983) );
  CMX2X1 U17204 ( .A0(n7971), .A1(n7983), .S(n4329), .Z(n7996) );
  CMXI2X1 U17205 ( .A0(n7972), .A1(n7996), .S(n3526), .Z(N2587) );
  CMX2X1 U17206 ( .A0(mem_data1[526]), .A1(mem_data1[527]), .S(n3878), .Z(
        n7979) );
  CMXI2X1 U17207 ( .A0(n7979), .A1(n7973), .S(n4042), .Z(n7986) );
  CMX2X1 U17208 ( .A0(n7974), .A1(n7986), .S(n4329), .Z(n8002) );
  CMXI2X1 U17209 ( .A0(n7975), .A1(n8002), .S(n3526), .Z(N2588) );
  CMX2X1 U17210 ( .A0(mem_data1[527]), .A1(mem_data1[528]), .S(n3879), .Z(
        n7982) );
  CMXI2X1 U17211 ( .A0(n7982), .A1(n7976), .S(n4042), .Z(n7989) );
  CMX2X1 U17212 ( .A0(n7977), .A1(n7989), .S(n4329), .Z(n8005) );
  CMXI2X1 U17213 ( .A0(n7978), .A1(n8005), .S(n3526), .Z(N2589) );
  CMX2X1 U17214 ( .A0(mem_data1[528]), .A1(mem_data1[529]), .S(n3869), .Z(
        n7985) );
  CMXI2X1 U17215 ( .A0(n7985), .A1(n7979), .S(n4042), .Z(n7992) );
  CMX2X1 U17216 ( .A0(n7980), .A1(n7992), .S(n4328), .Z(n8008) );
  CMXI2X1 U17217 ( .A0(n7981), .A1(n8008), .S(n3526), .Z(N2590) );
  CMX2X1 U17218 ( .A0(mem_data1[529]), .A1(mem_data1[530]), .S(n3870), .Z(
        n7988) );
  CMXI2X1 U17219 ( .A0(n7988), .A1(n7982), .S(n4042), .Z(n7995) );
  CMX2X1 U17220 ( .A0(n7983), .A1(n7995), .S(n4328), .Z(n8011) );
  CMXI2X1 U17221 ( .A0(n7984), .A1(n8011), .S(n3526), .Z(N2591) );
  CMX2X1 U17222 ( .A0(mem_data1[530]), .A1(mem_data1[531]), .S(n3871), .Z(
        n7991) );
  CMXI2X1 U17223 ( .A0(n7991), .A1(n7985), .S(n4042), .Z(n8001) );
  CMX2X1 U17224 ( .A0(n7986), .A1(n8001), .S(n4328), .Z(n8014) );
  CMXI2X1 U17225 ( .A0(n7987), .A1(n8014), .S(n3526), .Z(N2592) );
  CMX2X1 U17226 ( .A0(mem_data1[531]), .A1(mem_data1[532]), .S(n3872), .Z(
        n7994) );
  CMXI2X1 U17227 ( .A0(n7994), .A1(n7988), .S(n4042), .Z(n8004) );
  CMX2X1 U17228 ( .A0(n7989), .A1(n8004), .S(n4328), .Z(n8017) );
  CMXI2X1 U17229 ( .A0(n7990), .A1(n8017), .S(n3526), .Z(N2593) );
  CMX2X1 U17230 ( .A0(mem_data1[532]), .A1(mem_data1[533]), .S(n3870), .Z(
        n8000) );
  CMXI2X1 U17231 ( .A0(n8000), .A1(n7991), .S(n4042), .Z(n8007) );
  CMX2X1 U17232 ( .A0(n7992), .A1(n8007), .S(n4328), .Z(n8020) );
  CMXI2X1 U17233 ( .A0(n7993), .A1(n8020), .S(n3525), .Z(N2594) );
  CMX2X1 U17234 ( .A0(mem_data1[533]), .A1(mem_data1[534]), .S(n3862), .Z(
        n8003) );
  CMXI2X1 U17235 ( .A0(n8003), .A1(n7994), .S(n4042), .Z(n8010) );
  CMX2X1 U17236 ( .A0(n7995), .A1(n8010), .S(n4328), .Z(n8023) );
  CMXI2X1 U17237 ( .A0(n7996), .A1(n8023), .S(n3525), .Z(N2595) );
  CMX2X1 U17238 ( .A0(mem_data1[65]), .A1(mem_data1[66]), .S(n3863), .Z(n8063)
         );
  CMXI2X1 U17239 ( .A0(n8063), .A1(n7997), .S(n4042), .Z(n8130) );
  CMX2X1 U17240 ( .A0(n7998), .A1(n8130), .S(n4328), .Z(n8263) );
  CMXI2X1 U17241 ( .A0(n7999), .A1(n8263), .S(n3525), .Z(N2127) );
  CMX2X1 U17242 ( .A0(mem_data1[534]), .A1(mem_data1[535]), .S(n3864), .Z(
        n8006) );
  CMXI2X1 U17243 ( .A0(n8006), .A1(n8000), .S(n4041), .Z(n8013) );
  CMX2X1 U17244 ( .A0(n8001), .A1(n8013), .S(n4328), .Z(n8026) );
  CMXI2X1 U17245 ( .A0(n8002), .A1(n8026), .S(n3525), .Z(N2596) );
  CMX2X1 U17246 ( .A0(mem_data1[535]), .A1(mem_data1[536]), .S(n3865), .Z(
        n8009) );
  CMXI2X1 U17247 ( .A0(n8009), .A1(n8003), .S(n4041), .Z(n8016) );
  CMX2X1 U17248 ( .A0(n8004), .A1(n8016), .S(n4328), .Z(n8029) );
  CMXI2X1 U17249 ( .A0(n8005), .A1(n8029), .S(n3529), .Z(N2597) );
  CMX2X1 U17250 ( .A0(mem_data1[536]), .A1(mem_data1[537]), .S(n3866), .Z(
        n8012) );
  CMXI2X1 U17251 ( .A0(n8012), .A1(n8006), .S(n4041), .Z(n8019) );
  CMX2X1 U17252 ( .A0(n8007), .A1(n8019), .S(n4328), .Z(n8035) );
  CMXI2X1 U17253 ( .A0(n8008), .A1(n8035), .S(n3528), .Z(N2598) );
  CMX2X1 U17254 ( .A0(mem_data1[537]), .A1(mem_data1[538]), .S(n3867), .Z(
        n8015) );
  CMXI2X1 U17255 ( .A0(n8015), .A1(n8009), .S(n4041), .Z(n8022) );
  CMX2X1 U17256 ( .A0(n8010), .A1(n8022), .S(n4328), .Z(n8038) );
  CMXI2X1 U17257 ( .A0(n8011), .A1(n8038), .S(n3528), .Z(N2599) );
  CMX2X1 U17258 ( .A0(mem_data1[538]), .A1(mem_data1[539]), .S(n3868), .Z(
        n8018) );
  CMXI2X1 U17259 ( .A0(n8018), .A1(n8012), .S(n4041), .Z(n8025) );
  CMX2X1 U17260 ( .A0(n8013), .A1(n8025), .S(n4327), .Z(n8041) );
  CMXI2X1 U17261 ( .A0(n8014), .A1(n8041), .S(n3528), .Z(N2600) );
  CMX2X1 U17262 ( .A0(mem_data1[539]), .A1(mem_data1[540]), .S(n3880), .Z(
        n8021) );
  CMXI2X1 U17263 ( .A0(n8021), .A1(n8015), .S(n4041), .Z(n8028) );
  CMX2X1 U17264 ( .A0(n8016), .A1(n8028), .S(n4327), .Z(n8044) );
  CMXI2X1 U17265 ( .A0(n8017), .A1(n8044), .S(n3528), .Z(N2601) );
  CMX2X1 U17266 ( .A0(mem_data1[540]), .A1(mem_data1[541]), .S(n3881), .Z(
        n8024) );
  CMXI2X1 U17267 ( .A0(n8024), .A1(n8018), .S(n4041), .Z(n8034) );
  CMX2X1 U17268 ( .A0(n8019), .A1(n8034), .S(n4327), .Z(n8047) );
  CMXI2X1 U17269 ( .A0(n8020), .A1(n8047), .S(n3528), .Z(N2602) );
  CMX2X1 U17270 ( .A0(mem_data1[541]), .A1(mem_data1[542]), .S(n3869), .Z(
        n8027) );
  CMXI2X1 U17271 ( .A0(n8027), .A1(n8021), .S(n4041), .Z(n8037) );
  CMX2X1 U17272 ( .A0(n8022), .A1(n8037), .S(n4327), .Z(n8050) );
  CMXI2X1 U17273 ( .A0(n8023), .A1(n8050), .S(n3528), .Z(N2603) );
  CMX2X1 U17274 ( .A0(mem_data1[542]), .A1(mem_data1[543]), .S(n3870), .Z(
        n8033) );
  CMXI2X1 U17275 ( .A0(n8033), .A1(n8024), .S(n4041), .Z(n8040) );
  CMX2X1 U17276 ( .A0(n8025), .A1(n8040), .S(n4327), .Z(n8053) );
  CMXI2X1 U17277 ( .A0(n8026), .A1(n8053), .S(n3528), .Z(N2604) );
  CMX2X1 U17278 ( .A0(mem_data1[543]), .A1(mem_data1[544]), .S(n3880), .Z(
        n8036) );
  CMXI2X1 U17279 ( .A0(n8036), .A1(n8027), .S(n4041), .Z(n8043) );
  CMX2X1 U17280 ( .A0(n8028), .A1(n8043), .S(n4327), .Z(n8056) );
  CMXI2X1 U17281 ( .A0(n8029), .A1(n8056), .S(n3528), .Z(N2605) );
  CMX2X1 U17282 ( .A0(mem_data1[66]), .A1(mem_data1[67]), .S(n3881), .Z(n8096)
         );
  CMXI2X1 U17283 ( .A0(n8096), .A1(n8030), .S(n4041), .Z(n8163) );
  CMX2X1 U17284 ( .A0(n8031), .A1(n8163), .S(n4327), .Z(n8300) );
  CMXI2X1 U17285 ( .A0(n8032), .A1(n8300), .S(n3527), .Z(N2128) );
  CMX2X1 U17286 ( .A0(mem_data1[544]), .A1(mem_data1[545]), .S(n3862), .Z(
        n8039) );
  CMXI2X1 U17287 ( .A0(n8039), .A1(n8033), .S(n4041), .Z(n8046) );
  CMX2X1 U17288 ( .A0(n8034), .A1(n8046), .S(n4327), .Z(n8059) );
  CMXI2X1 U17289 ( .A0(n8035), .A1(n8059), .S(n3528), .Z(N2606) );
  CMX2X1 U17290 ( .A0(mem_data1[545]), .A1(mem_data1[546]), .S(n3863), .Z(
        n8042) );
  CMXI2X1 U17291 ( .A0(n8042), .A1(n8036), .S(n4041), .Z(n8049) );
  CMX2X1 U17292 ( .A0(n8037), .A1(n8049), .S(n4327), .Z(n8062) );
  CMXI2X1 U17293 ( .A0(n8038), .A1(n8062), .S(n3527), .Z(N2607) );
  CMX2X1 U17294 ( .A0(mem_data1[546]), .A1(mem_data1[547]), .S(n3873), .Z(
        n8045) );
  CMXI2X1 U17295 ( .A0(n8045), .A1(n8039), .S(n4041), .Z(n8052) );
  CMX2X1 U17296 ( .A0(n8040), .A1(n8052), .S(n4327), .Z(n8068) );
  CMXI2X1 U17297 ( .A0(n8041), .A1(n8068), .S(n3527), .Z(N2608) );
  CMX2X1 U17298 ( .A0(mem_data1[547]), .A1(mem_data1[548]), .S(n3874), .Z(
        n8048) );
  CMXI2X1 U17299 ( .A0(n8048), .A1(n8042), .S(n4041), .Z(n8055) );
  CMX2X1 U17300 ( .A0(n8043), .A1(n8055), .S(n4327), .Z(n8071) );
  CMXI2X1 U17301 ( .A0(n8044), .A1(n8071), .S(n3527), .Z(N2609) );
  CMX2X1 U17302 ( .A0(mem_data1[548]), .A1(mem_data1[549]), .S(n3875), .Z(
        n8051) );
  CMXI2X1 U17303 ( .A0(n8051), .A1(n8045), .S(n4041), .Z(n8058) );
  CMX2X1 U17304 ( .A0(n8046), .A1(n8058), .S(n4326), .Z(n8074) );
  CMXI2X1 U17305 ( .A0(n8047), .A1(n8074), .S(n3527), .Z(N2610) );
  CMX2X1 U17306 ( .A0(mem_data1[549]), .A1(mem_data1[550]), .S(n3876), .Z(
        n8054) );
  CMXI2X1 U17307 ( .A0(n8054), .A1(n8048), .S(n4040), .Z(n8061) );
  CMX2X1 U17308 ( .A0(n8049), .A1(n8061), .S(n4326), .Z(n8077) );
  CMXI2X1 U17309 ( .A0(n8050), .A1(n8077), .S(n3527), .Z(N2611) );
  CMX2X1 U17310 ( .A0(mem_data1[550]), .A1(mem_data1[551]), .S(n3871), .Z(
        n8057) );
  CMXI2X1 U17311 ( .A0(n8057), .A1(n8051), .S(n4040), .Z(n8067) );
  CMX2X1 U17312 ( .A0(n8052), .A1(n8067), .S(n4326), .Z(n8080) );
  CMXI2X1 U17313 ( .A0(n8053), .A1(n8080), .S(n3527), .Z(N2612) );
  CMX2X1 U17314 ( .A0(mem_data1[551]), .A1(mem_data1[552]), .S(n3871), .Z(
        n8060) );
  CMXI2X1 U17315 ( .A0(n8060), .A1(n8054), .S(n4040), .Z(n8070) );
  CMX2X1 U17316 ( .A0(n8055), .A1(n8070), .S(n4326), .Z(n8083) );
  CMXI2X1 U17317 ( .A0(n8056), .A1(n8083), .S(n3527), .Z(N2613) );
  CMX2X1 U17318 ( .A0(mem_data1[552]), .A1(mem_data1[553]), .S(n3872), .Z(
        n8066) );
  CMXI2X1 U17319 ( .A0(n8066), .A1(n8057), .S(n4040), .Z(n8073) );
  CMX2X1 U17320 ( .A0(n8058), .A1(n8073), .S(n4326), .Z(n8086) );
  CMXI2X1 U17321 ( .A0(n8059), .A1(n8086), .S(n3529), .Z(N2614) );
  CMX2X1 U17322 ( .A0(mem_data1[553]), .A1(mem_data1[554]), .S(n3873), .Z(
        n8069) );
  CMXI2X1 U17323 ( .A0(n8069), .A1(n8060), .S(n4040), .Z(n8076) );
  CMX2X1 U17324 ( .A0(n8061), .A1(n8076), .S(n4326), .Z(n8089) );
  CMXI2X1 U17325 ( .A0(n8062), .A1(n8089), .S(n3530), .Z(N2615) );
  CMX2X1 U17326 ( .A0(mem_data1[67]), .A1(mem_data1[68]), .S(n3874), .Z(n8129)
         );
  CMXI2X1 U17327 ( .A0(n8129), .A1(n8063), .S(n4040), .Z(n8196) );
  CMX2X1 U17328 ( .A0(n8064), .A1(n8196), .S(n4326), .Z(n8333) );
  CMXI2X1 U17329 ( .A0(n8065), .A1(n8333), .S(n3530), .Z(N2129) );
  CMX2X1 U17330 ( .A0(mem_data1[554]), .A1(mem_data1[555]), .S(n3875), .Z(
        n8072) );
  CMXI2X1 U17331 ( .A0(n8072), .A1(n8066), .S(n4040), .Z(n8079) );
  CMX2X1 U17332 ( .A0(n8067), .A1(n8079), .S(n4326), .Z(n8092) );
  CMXI2X1 U17333 ( .A0(n8068), .A1(n8092), .S(n3530), .Z(N2616) );
  CMX2X1 U17334 ( .A0(mem_data1[555]), .A1(mem_data1[556]), .S(n3876), .Z(
        n8075) );
  CMXI2X1 U17335 ( .A0(n8075), .A1(n8069), .S(n4040), .Z(n8082) );
  CMX2X1 U17336 ( .A0(n8070), .A1(n8082), .S(n4326), .Z(n8095) );
  CMXI2X1 U17337 ( .A0(n8071), .A1(n8095), .S(n3529), .Z(N2617) );
  CMX2X1 U17338 ( .A0(mem_data1[556]), .A1(mem_data1[557]), .S(n3877), .Z(
        n8078) );
  CMXI2X1 U17339 ( .A0(n8078), .A1(n8072), .S(n4040), .Z(n8085) );
  CMX2X1 U17340 ( .A0(n8073), .A1(n8085), .S(n4326), .Z(n8101) );
  CMXI2X1 U17341 ( .A0(n8074), .A1(n8101), .S(n3530), .Z(N2618) );
  CMX2X1 U17342 ( .A0(mem_data1[557]), .A1(mem_data1[558]), .S(n3862), .Z(
        n8081) );
  CMXI2X1 U17343 ( .A0(n8081), .A1(n8075), .S(n4040), .Z(n8088) );
  CMX2X1 U17344 ( .A0(n8076), .A1(n8088), .S(n4326), .Z(n8104) );
  CMXI2X1 U17345 ( .A0(n8077), .A1(n8104), .S(n3530), .Z(N2619) );
  CMX2X1 U17346 ( .A0(mem_data1[558]), .A1(mem_data1[559]), .S(n3863), .Z(
        n8084) );
  CMXI2X1 U17347 ( .A0(n8084), .A1(n8078), .S(n4040), .Z(n8091) );
  CMX2X1 U17348 ( .A0(n8079), .A1(n8091), .S(n4325), .Z(n8107) );
  CMXI2X1 U17349 ( .A0(n8080), .A1(n8107), .S(n3530), .Z(N2620) );
  CMX2X1 U17350 ( .A0(mem_data1[559]), .A1(mem_data1[560]), .S(n3878), .Z(
        n8087) );
  CMXI2X1 U17351 ( .A0(n8087), .A1(n8081), .S(n4040), .Z(n8094) );
  CMX2X1 U17352 ( .A0(n8082), .A1(n8094), .S(n4325), .Z(n8110) );
  CMXI2X1 U17353 ( .A0(n8083), .A1(n8110), .S(n3529), .Z(N2621) );
  CMX2X1 U17354 ( .A0(mem_data1[560]), .A1(mem_data1[561]), .S(n3879), .Z(
        n8090) );
  CMXI2X1 U17355 ( .A0(n8090), .A1(n8084), .S(n4040), .Z(n8100) );
  CMX2X1 U17356 ( .A0(n8085), .A1(n8100), .S(n4325), .Z(n8113) );
  CMXI2X1 U17357 ( .A0(n8086), .A1(n8113), .S(n3529), .Z(N2622) );
  CMX2X1 U17358 ( .A0(mem_data1[561]), .A1(mem_data1[562]), .S(n3864), .Z(
        n8093) );
  CMXI2X1 U17359 ( .A0(n8093), .A1(n8087), .S(n4040), .Z(n8103) );
  CMX2X1 U17360 ( .A0(n8088), .A1(n8103), .S(n4325), .Z(n8116) );
  CMXI2X1 U17361 ( .A0(n8089), .A1(n8116), .S(n3529), .Z(N2623) );
  CMX2X1 U17362 ( .A0(mem_data1[562]), .A1(mem_data1[563]), .S(n3865), .Z(
        n8099) );
  CMXI2X1 U17363 ( .A0(n8099), .A1(n8090), .S(n4040), .Z(n8106) );
  CMX2X1 U17364 ( .A0(n8091), .A1(n8106), .S(n4325), .Z(n8119) );
  CMXI2X1 U17365 ( .A0(n8092), .A1(n8119), .S(n3529), .Z(N2624) );
  CMX2X1 U17366 ( .A0(mem_data1[563]), .A1(mem_data1[564]), .S(n3866), .Z(
        n8102) );
  CMXI2X1 U17367 ( .A0(n8102), .A1(n8093), .S(n4040), .Z(n8109) );
  CMX2X1 U17368 ( .A0(n8094), .A1(n8109), .S(n4325), .Z(n8122) );
  CMXI2X1 U17369 ( .A0(n8095), .A1(n8122), .S(n3528), .Z(N2625) );
  CMX2X1 U17370 ( .A0(mem_data1[68]), .A1(mem_data1[69]), .S(n3867), .Z(n8162)
         );
  CMXI2X1 U17371 ( .A0(n8162), .A1(n8096), .S(n4039), .Z(n8229) );
  CMX2X1 U17372 ( .A0(n8097), .A1(n8229), .S(n4325), .Z(n8366) );
  CMXI2X1 U17373 ( .A0(n8098), .A1(n8366), .S(n3529), .Z(N2130) );
  CMX2X1 U17374 ( .A0(mem_data1[564]), .A1(mem_data1[565]), .S(n3877), .Z(
        n8105) );
  CMXI2X1 U17375 ( .A0(n8105), .A1(n8099), .S(n4039), .Z(n8112) );
  CMX2X1 U17376 ( .A0(n8100), .A1(n8112), .S(n4325), .Z(n8125) );
  CMXI2X1 U17377 ( .A0(n8101), .A1(n8125), .S(n3529), .Z(N2626) );
  CMX2X1 U17378 ( .A0(mem_data1[565]), .A1(mem_data1[566]), .S(n3878), .Z(
        n8108) );
  CMXI2X1 U17379 ( .A0(n8108), .A1(n8102), .S(n4039), .Z(n8115) );
  CMX2X1 U17380 ( .A0(n8103), .A1(n8115), .S(n4325), .Z(n8128) );
  CMXI2X1 U17381 ( .A0(n8104), .A1(n8128), .S(n3529), .Z(N2627) );
  CMX2X1 U17382 ( .A0(mem_data1[566]), .A1(mem_data1[567]), .S(n3879), .Z(
        n8111) );
  CMXI2X1 U17383 ( .A0(n8111), .A1(n8105), .S(n4039), .Z(n8118) );
  CMX2X1 U17384 ( .A0(n8106), .A1(n8118), .S(n4325), .Z(n8134) );
  CMXI2X1 U17385 ( .A0(n8107), .A1(n8134), .S(n3528), .Z(N2628) );
  CMX2X1 U17386 ( .A0(mem_data1[567]), .A1(mem_data1[568]), .S(n3880), .Z(
        n8114) );
  CMXI2X1 U17387 ( .A0(n8114), .A1(n8108), .S(n4039), .Z(n8121) );
  CMX2X1 U17388 ( .A0(n8109), .A1(n8121), .S(n4325), .Z(n8137) );
  CMXI2X1 U17389 ( .A0(n8110), .A1(n8137), .S(n3529), .Z(N2629) );
  CMX2X1 U17390 ( .A0(mem_data1[568]), .A1(mem_data1[569]), .S(n3872), .Z(
        n8117) );
  CMXI2X1 U17391 ( .A0(n8117), .A1(n8111), .S(n4039), .Z(n8124) );
  CMX2X1 U17392 ( .A0(n8112), .A1(n8124), .S(n4324), .Z(n8140) );
  CMXI2X1 U17393 ( .A0(n8113), .A1(n8140), .S(n3532), .Z(N2630) );
  CMX2X1 U17394 ( .A0(mem_data1[569]), .A1(mem_data1[570]), .S(n3880), .Z(
        n8120) );
  CMXI2X1 U17395 ( .A0(n8120), .A1(n8114), .S(n4039), .Z(n8127) );
  CMX2X1 U17396 ( .A0(n8115), .A1(n8127), .S(n4324), .Z(n8143) );
  CMXI2X1 U17397 ( .A0(n8116), .A1(n8143), .S(n3532), .Z(N2631) );
  CMX2X1 U17398 ( .A0(mem_data1[570]), .A1(mem_data1[571]), .S(n3881), .Z(
        n8123) );
  CMXI2X1 U17399 ( .A0(n8123), .A1(n8117), .S(n4039), .Z(n8133) );
  CMX2X1 U17400 ( .A0(n8118), .A1(n8133), .S(n4324), .Z(n8146) );
  CMXI2X1 U17401 ( .A0(n8119), .A1(n8146), .S(n3531), .Z(N2632) );
  CMX2X1 U17402 ( .A0(mem_data1[571]), .A1(mem_data1[572]), .S(n3862), .Z(
        n8126) );
  CMXI2X1 U17403 ( .A0(n8126), .A1(n8120), .S(n4039), .Z(n8136) );
  CMX2X1 U17404 ( .A0(n8121), .A1(n8136), .S(n4324), .Z(n8149) );
  CMXI2X1 U17405 ( .A0(n8122), .A1(n8149), .S(n3532), .Z(N2633) );
  CMX2X1 U17406 ( .A0(mem_data1[572]), .A1(mem_data1[573]), .S(n3863), .Z(
        n8132) );
  CMXI2X1 U17407 ( .A0(n8132), .A1(n8123), .S(n4039), .Z(n8139) );
  CMX2X1 U17408 ( .A0(n8124), .A1(n8139), .S(n4324), .Z(n8152) );
  CMXI2X1 U17409 ( .A0(n8125), .A1(n8152), .S(n3531), .Z(N2634) );
  CMX2X1 U17410 ( .A0(mem_data1[573]), .A1(mem_data1[574]), .S(n3864), .Z(
        n8135) );
  CMXI2X1 U17411 ( .A0(n8135), .A1(n8126), .S(n4039), .Z(n8142) );
  CMX2X1 U17412 ( .A0(n8127), .A1(n8142), .S(n4324), .Z(n8155) );
  CMXI2X1 U17413 ( .A0(n8128), .A1(n8155), .S(n3531), .Z(N2635) );
  CMX2X1 U17414 ( .A0(mem_data1[69]), .A1(mem_data1[70]), .S(n3865), .Z(n8195)
         );
  CMXI2X1 U17415 ( .A0(n8195), .A1(n8129), .S(n4039), .Z(n8262) );
  CMX2X1 U17416 ( .A0(n8130), .A1(n8262), .S(n4324), .Z(n8399) );
  CMXI2X1 U17417 ( .A0(n8131), .A1(n8399), .S(n3531), .Z(N2131) );
  CMX2X1 U17418 ( .A0(mem_data1[574]), .A1(mem_data1[575]), .S(n3866), .Z(
        n8138) );
  CMXI2X1 U17419 ( .A0(n8138), .A1(n8132), .S(n4039), .Z(n8145) );
  CMX2X1 U17420 ( .A0(n8133), .A1(n8145), .S(n4324), .Z(n8158) );
  CMXI2X1 U17421 ( .A0(n8134), .A1(n8158), .S(n3531), .Z(N2636) );
  CMX2X1 U17422 ( .A0(mem_data1[575]), .A1(mem_data1[576]), .S(n3864), .Z(
        n8141) );
  CMXI2X1 U17423 ( .A0(n8141), .A1(n8135), .S(n4039), .Z(n8148) );
  CMX2X1 U17424 ( .A0(n8136), .A1(n8148), .S(n4324), .Z(n8161) );
  CMXI2X1 U17425 ( .A0(n8137), .A1(n8161), .S(n3531), .Z(N2637) );
  CMX2X1 U17426 ( .A0(mem_data1[576]), .A1(mem_data1[577]), .S(n3865), .Z(
        n8144) );
  CMXI2X1 U17427 ( .A0(n8144), .A1(n8138), .S(n4039), .Z(n8151) );
  CMX2X1 U17428 ( .A0(n8139), .A1(n8151), .S(n4324), .Z(n8167) );
  CMXI2X1 U17429 ( .A0(n8140), .A1(n8167), .S(n3531), .Z(N2638) );
  CMX2X1 U17430 ( .A0(mem_data1[577]), .A1(mem_data1[578]), .S(n3867), .Z(
        n8147) );
  CMXI2X1 U17431 ( .A0(n8147), .A1(n8141), .S(n4039), .Z(n8154) );
  CMX2X1 U17432 ( .A0(n8142), .A1(n8154), .S(n4324), .Z(n8170) );
  CMXI2X1 U17433 ( .A0(n8143), .A1(n8170), .S(n3530), .Z(N2639) );
  CMX2X1 U17434 ( .A0(mem_data1[578]), .A1(mem_data1[579]), .S(n3868), .Z(
        n8150) );
  CMXI2X1 U17435 ( .A0(n8150), .A1(n8144), .S(n4038), .Z(n8157) );
  CMX2X1 U17436 ( .A0(n8145), .A1(n8157), .S(n4323), .Z(n8173) );
  CMXI2X1 U17437 ( .A0(n8146), .A1(n8173), .S(n3531), .Z(N2640) );
  CMX2X1 U17438 ( .A0(mem_data1[579]), .A1(mem_data1[580]), .S(n3868), .Z(
        n8153) );
  CMXI2X1 U17439 ( .A0(n8153), .A1(n8147), .S(n4038), .Z(n8160) );
  CMX2X1 U17440 ( .A0(n8148), .A1(n8160), .S(n4323), .Z(n8176) );
  CMXI2X1 U17441 ( .A0(n8149), .A1(n8176), .S(n3531), .Z(N2641) );
  CMX2X1 U17442 ( .A0(mem_data1[580]), .A1(mem_data1[581]), .S(n3869), .Z(
        n8156) );
  CMXI2X1 U17443 ( .A0(n8156), .A1(n8150), .S(n4038), .Z(n8166) );
  CMX2X1 U17444 ( .A0(n8151), .A1(n8166), .S(n4323), .Z(n8179) );
  CMXI2X1 U17445 ( .A0(n8152), .A1(n8179), .S(n3531), .Z(N2642) );
  CMX2X1 U17446 ( .A0(mem_data1[581]), .A1(mem_data1[582]), .S(n3870), .Z(
        n8159) );
  CMXI2X1 U17447 ( .A0(n8159), .A1(n8153), .S(n4038), .Z(n8169) );
  CMX2X1 U17448 ( .A0(n8154), .A1(n8169), .S(n4323), .Z(n8182) );
  CMXI2X1 U17449 ( .A0(n8155), .A1(n8182), .S(n3530), .Z(N2643) );
  CMX2X1 U17450 ( .A0(mem_data1[582]), .A1(mem_data1[583]), .S(n3871), .Z(
        n8165) );
  CMXI2X1 U17451 ( .A0(n8165), .A1(n8156), .S(n4038), .Z(n8172) );
  CMX2X1 U17452 ( .A0(n8157), .A1(n8172), .S(n4323), .Z(n8185) );
  CMXI2X1 U17453 ( .A0(n8158), .A1(n8185), .S(n3530), .Z(N2644) );
  CMX2X1 U17454 ( .A0(mem_data1[583]), .A1(mem_data1[584]), .S(n3881), .Z(
        n8168) );
  CMXI2X1 U17455 ( .A0(n8168), .A1(n8159), .S(n4038), .Z(n8175) );
  CMX2X1 U17456 ( .A0(n8160), .A1(n8175), .S(n4323), .Z(n8188) );
  CMXI2X1 U17457 ( .A0(n8161), .A1(n8188), .S(n3530), .Z(N2645) );
  CMX2X1 U17458 ( .A0(mem_data1[70]), .A1(mem_data1[71]), .S(n3862), .Z(n8228)
         );
  CMXI2X1 U17459 ( .A0(n8228), .A1(n8162), .S(n4038), .Z(n8299) );
  CMX2X1 U17460 ( .A0(n8163), .A1(n8299), .S(n4323), .Z(n8432) );
  CMXI2X1 U17461 ( .A0(n8164), .A1(n8432), .S(n3530), .Z(N2132) );
  CMX2X1 U17462 ( .A0(mem_data1[584]), .A1(mem_data1[585]), .S(n3863), .Z(
        n8171) );
  CMXI2X1 U17463 ( .A0(n8171), .A1(n8165), .S(n4038), .Z(n8178) );
  CMX2X1 U17464 ( .A0(n8166), .A1(n8178), .S(n4323), .Z(n8191) );
  CMXI2X1 U17465 ( .A0(n8167), .A1(n8191), .S(n3499), .Z(N2646) );
  CMX2X1 U17466 ( .A0(mem_data1[585]), .A1(mem_data1[586]), .S(n3878), .Z(
        n8174) );
  CMXI2X1 U17467 ( .A0(n8174), .A1(n8168), .S(n4038), .Z(n8181) );
  CMX2X1 U17468 ( .A0(n8169), .A1(n8181), .S(n4323), .Z(n8194) );
  CMXI2X1 U17469 ( .A0(n8170), .A1(n8194), .S(n3499), .Z(N2647) );
  CMX2X1 U17470 ( .A0(mem_data1[586]), .A1(mem_data1[587]), .S(n3870), .Z(
        n8177) );
  CMXI2X1 U17471 ( .A0(n8177), .A1(n8171), .S(n4038), .Z(n8184) );
  CMX2X1 U17472 ( .A0(n8172), .A1(n8184), .S(n4323), .Z(n8200) );
  CMXI2X1 U17473 ( .A0(n8173), .A1(n8200), .S(n3499), .Z(N2648) );
  CMX2X1 U17474 ( .A0(mem_data1[587]), .A1(mem_data1[588]), .S(n3871), .Z(
        n8180) );
  CMXI2X1 U17475 ( .A0(n8180), .A1(n8174), .S(n4038), .Z(n8187) );
  CMX2X1 U17476 ( .A0(n8175), .A1(n8187), .S(n4323), .Z(n8203) );
  CMXI2X1 U17477 ( .A0(n8176), .A1(n8203), .S(n3498), .Z(N2649) );
  CMX2X1 U17478 ( .A0(mem_data1[588]), .A1(mem_data1[589]), .S(n3874), .Z(
        n8183) );
  CMXI2X1 U17479 ( .A0(n8183), .A1(n8177), .S(n4038), .Z(n8190) );
  CMX2X1 U17480 ( .A0(n8178), .A1(n8190), .S(n4322), .Z(n8206) );
  CMXI2X1 U17481 ( .A0(n8179), .A1(n8206), .S(n3498), .Z(N2650) );
  CMX2X1 U17482 ( .A0(mem_data1[589]), .A1(mem_data1[590]), .S(n3864), .Z(
        n8186) );
  CMXI2X1 U17483 ( .A0(n8186), .A1(n8180), .S(n4038), .Z(n8193) );
  CMX2X1 U17484 ( .A0(n8181), .A1(n8193), .S(n4322), .Z(n8209) );
  CMXI2X1 U17485 ( .A0(n8182), .A1(n8209), .S(n3498), .Z(N2651) );
  CMX2X1 U17486 ( .A0(mem_data1[590]), .A1(mem_data1[591]), .S(n3865), .Z(
        n8189) );
  CMXI2X1 U17487 ( .A0(n8189), .A1(n8183), .S(n4038), .Z(n8199) );
  CMX2X1 U17488 ( .A0(n8184), .A1(n8199), .S(n4322), .Z(n8212) );
  CMXI2X1 U17489 ( .A0(n8185), .A1(n8212), .S(n3498), .Z(N2652) );
  CMX2X1 U17490 ( .A0(mem_data1[591]), .A1(mem_data1[592]), .S(n3866), .Z(
        n8192) );
  CMXI2X1 U17491 ( .A0(n8192), .A1(n8186), .S(n4038), .Z(n8202) );
  CMX2X1 U17492 ( .A0(n8187), .A1(n8202), .S(n4322), .Z(n8215) );
  CMXI2X1 U17493 ( .A0(n8188), .A1(n8215), .S(n3498), .Z(N2653) );
  CMX2X1 U17494 ( .A0(mem_data1[592]), .A1(mem_data1[593]), .S(n3867), .Z(
        n8198) );
  CMXI2X1 U17495 ( .A0(n8198), .A1(n8189), .S(n4038), .Z(n8205) );
  CMX2X1 U17496 ( .A0(n8190), .A1(n8205), .S(n4322), .Z(n8218) );
  CMXI2X1 U17497 ( .A0(n8191), .A1(n8218), .S(n3498), .Z(N2654) );
  CMX2X1 U17498 ( .A0(mem_data1[593]), .A1(mem_data1[594]), .S(n3868), .Z(
        n8201) );
  CMXI2X1 U17499 ( .A0(n8201), .A1(n8192), .S(n4037), .Z(n8208) );
  CMX2X1 U17500 ( .A0(n8193), .A1(n8208), .S(n4322), .Z(n8221) );
  CMXI2X1 U17501 ( .A0(n8194), .A1(n8221), .S(n3507), .Z(N2655) );
  CMX2X1 U17502 ( .A0(mem_data1[71]), .A1(mem_data1[72]), .S(n3869), .Z(n8261)
         );
  CMXI2X1 U17503 ( .A0(n8261), .A1(n8195), .S(n4037), .Z(n8332) );
  CMX2X1 U17504 ( .A0(n8196), .A1(n8332), .S(n4322), .Z(n8465) );
  CMXI2X1 U17505 ( .A0(n8197), .A1(n8465), .S(n3532), .Z(N2133) );
  CMX2X1 U17506 ( .A0(mem_data1[594]), .A1(mem_data1[595]), .S(n3870), .Z(
        n8204) );
  CMXI2X1 U17507 ( .A0(n8204), .A1(n8198), .S(n4037), .Z(n8211) );
  CMX2X1 U17508 ( .A0(n8199), .A1(n8211), .S(n4322), .Z(n8224) );
  CMXI2X1 U17509 ( .A0(n8200), .A1(n8224), .S(n3532), .Z(N2656) );
  CMX2X1 U17510 ( .A0(mem_data1[595]), .A1(mem_data1[596]), .S(n3880), .Z(
        n8207) );
  CMXI2X1 U17511 ( .A0(n8207), .A1(n8201), .S(n4037), .Z(n8214) );
  CMX2X1 U17512 ( .A0(n8202), .A1(n8214), .S(n4322), .Z(n8227) );
  CMXI2X1 U17513 ( .A0(n8203), .A1(n8227), .S(n3532), .Z(N2657) );
  CMX2X1 U17514 ( .A0(mem_data1[596]), .A1(mem_data1[597]), .S(n3881), .Z(
        n8210) );
  CMXI2X1 U17515 ( .A0(n8210), .A1(n8204), .S(n4037), .Z(n8217) );
  CMX2X1 U17516 ( .A0(n8205), .A1(n8217), .S(n4330), .Z(n8233) );
  CMXI2X1 U17517 ( .A0(n8206), .A1(n8233), .S(n3532), .Z(N2658) );
  CMX2X1 U17518 ( .A0(mem_data1[597]), .A1(mem_data1[598]), .S(n3871), .Z(
        n8213) );
  CMXI2X1 U17519 ( .A0(n8213), .A1(n8207), .S(n4037), .Z(n8220) );
  CMX2X1 U17520 ( .A0(n8208), .A1(n8220), .S(n4353), .Z(n8236) );
  CMXI2X1 U17521 ( .A0(n8209), .A1(n8236), .S(n3532), .Z(N2659) );
  CMX2X1 U17522 ( .A0(mem_data1[598]), .A1(mem_data1[599]), .S(n3872), .Z(
        n8216) );
  CMXI2X1 U17523 ( .A0(n8216), .A1(n8210), .S(n4037), .Z(n8223) );
  CMX2X1 U17524 ( .A0(n8211), .A1(n8223), .S(n4353), .Z(n8239) );
  CMXI2X1 U17525 ( .A0(n8212), .A1(n8239), .S(n3532), .Z(N2660) );
  CMX2X1 U17526 ( .A0(mem_data1[599]), .A1(mem_data1[600]), .S(n3864), .Z(
        n8219) );
  CMXI2X1 U17527 ( .A0(n8219), .A1(n8213), .S(n4037), .Z(n8226) );
  CMX2X1 U17528 ( .A0(n8214), .A1(n8226), .S(n4353), .Z(n8242) );
  CMXI2X1 U17529 ( .A0(n8215), .A1(n8242), .S(n3531), .Z(N2661) );
  CMX2X1 U17530 ( .A0(mem_data1[600]), .A1(mem_data1[601]), .S(n3865), .Z(
        n8222) );
  CMXI2X1 U17531 ( .A0(n8222), .A1(n8216), .S(n4037), .Z(n8232) );
  CMX2X1 U17532 ( .A0(n8217), .A1(n8232), .S(n4353), .Z(n8245) );
  CMXI2X1 U17533 ( .A0(n8218), .A1(n8245), .S(n3532), .Z(N2662) );
  CMX2X1 U17534 ( .A0(mem_data1[601]), .A1(mem_data1[602]), .S(n3866), .Z(
        n8225) );
  CMXI2X1 U17535 ( .A0(n8225), .A1(n8219), .S(n4037), .Z(n8235) );
  CMX2X1 U17536 ( .A0(n8220), .A1(n8235), .S(n4353), .Z(n8248) );
  CMXI2X1 U17537 ( .A0(n8221), .A1(n8248), .S(n3350), .Z(N2663) );
  CMX2X1 U17538 ( .A0(mem_data1[602]), .A1(mem_data1[603]), .S(n3867), .Z(
        n8231) );
  CMXI2X1 U17539 ( .A0(n8231), .A1(n8222), .S(n4037), .Z(n8238) );
  CMX2X1 U17540 ( .A0(n8223), .A1(n8238), .S(n4353), .Z(n8251) );
  CMXI2X1 U17541 ( .A0(n8224), .A1(n8251), .S(n3350), .Z(N2664) );
  CMX2X1 U17542 ( .A0(mem_data1[603]), .A1(mem_data1[604]), .S(n3864), .Z(
        n8234) );
  CMXI2X1 U17543 ( .A0(n8234), .A1(n8225), .S(n4037), .Z(n8241) );
  CMX2X1 U17544 ( .A0(n8226), .A1(n8241), .S(n4352), .Z(n8254) );
  CMXI2X1 U17545 ( .A0(n8227), .A1(n8254), .S(n3350), .Z(N2665) );
  CMX2X1 U17546 ( .A0(mem_data1[72]), .A1(mem_data1[73]), .S(n3865), .Z(n8298)
         );
  CMXI2X1 U17547 ( .A0(n8298), .A1(n8228), .S(n4037), .Z(n8365) );
  CMX2X1 U17548 ( .A0(n8229), .A1(n8365), .S(n4352), .Z(n8498) );
  CMXI2X1 U17549 ( .A0(n8230), .A1(n8498), .S(n3350), .Z(N2134) );
  CMX2X1 U17550 ( .A0(mem_data1[604]), .A1(mem_data1[605]), .S(n3866), .Z(
        n8237) );
  CMXI2X1 U17551 ( .A0(n8237), .A1(n8231), .S(n4037), .Z(n8244) );
  CMX2X1 U17552 ( .A0(n8232), .A1(n8244), .S(n4352), .Z(n8257) );
  CMXI2X1 U17553 ( .A0(n8233), .A1(n8257), .S(n3349), .Z(N2666) );
  CMX2X1 U17554 ( .A0(mem_data1[605]), .A1(mem_data1[606]), .S(n3867), .Z(
        n8240) );
  CMXI2X1 U17555 ( .A0(n8240), .A1(n8234), .S(n4037), .Z(n8247) );
  CMX2X1 U17556 ( .A0(n8235), .A1(n8247), .S(n4352), .Z(n8260) );
  CMXI2X1 U17557 ( .A0(n8236), .A1(n8260), .S(n3349), .Z(N2667) );
  CMX2X1 U17558 ( .A0(mem_data1[606]), .A1(mem_data1[607]), .S(n3872), .Z(
        n8243) );
  CMXI2X1 U17559 ( .A0(n8243), .A1(n8237), .S(n4037), .Z(n8250) );
  CMX2X1 U17560 ( .A0(n8238), .A1(n8250), .S(n4352), .Z(n8270) );
  CMXI2X1 U17561 ( .A0(n8239), .A1(n8270), .S(n3349), .Z(N2668) );
  CMX2X1 U17562 ( .A0(mem_data1[607]), .A1(mem_data1[608]), .S(n3873), .Z(
        n8246) );
  CMXI2X1 U17563 ( .A0(n8246), .A1(n8240), .S(n4036), .Z(n8253) );
  CMX2X1 U17564 ( .A0(n8241), .A1(n8253), .S(n4352), .Z(n8273) );
  CMXI2X1 U17565 ( .A0(n8242), .A1(n8273), .S(n3349), .Z(N2669) );
  CMX2X1 U17566 ( .A0(mem_data1[608]), .A1(mem_data1[609]), .S(n3874), .Z(
        n8249) );
  CMXI2X1 U17567 ( .A0(n8249), .A1(n8243), .S(n4036), .Z(n8256) );
  CMX2X1 U17568 ( .A0(n8244), .A1(n8256), .S(n4352), .Z(n8276) );
  CMXI2X1 U17569 ( .A0(n8245), .A1(n8276), .S(n3349), .Z(N2670) );
  CMX2X1 U17570 ( .A0(mem_data1[609]), .A1(mem_data1[610]), .S(n3875), .Z(
        n8252) );
  CMXI2X1 U17571 ( .A0(n8252), .A1(n8246), .S(n4036), .Z(n8259) );
  CMX2X1 U17572 ( .A0(n8247), .A1(n8259), .S(n4352), .Z(n8279) );
  CMXI2X1 U17573 ( .A0(n8248), .A1(n8279), .S(n3349), .Z(N2671) );
  CMX2X1 U17574 ( .A0(mem_data1[610]), .A1(mem_data1[611]), .S(n3872), .Z(
        n8255) );
  CMXI2X1 U17575 ( .A0(n8255), .A1(n8249), .S(n4036), .Z(n8269) );
  CMX2X1 U17576 ( .A0(n8250), .A1(n8269), .S(n4352), .Z(n8282) );
  CMXI2X1 U17577 ( .A0(n8251), .A1(n8282), .S(n3349), .Z(N2672) );
  CMX2X1 U17578 ( .A0(mem_data1[611]), .A1(mem_data1[612]), .S(n3873), .Z(
        n8258) );
  CMXI2X1 U17579 ( .A0(n8258), .A1(n8252), .S(n4036), .Z(n8272) );
  CMX2X1 U17580 ( .A0(n8253), .A1(n8272), .S(n4352), .Z(n8285) );
  CMXI2X1 U17581 ( .A0(n8254), .A1(n8285), .S(n3473), .Z(N2673) );
  CMX2X1 U17582 ( .A0(mem_data1[612]), .A1(mem_data1[613]), .S(n3868), .Z(
        n8268) );
  CMXI2X1 U17583 ( .A0(n8268), .A1(n8255), .S(n4036), .Z(n8275) );
  CMX2X1 U17584 ( .A0(n8256), .A1(n8275), .S(n4352), .Z(n8288) );
  CMXI2X1 U17585 ( .A0(n8257), .A1(n8288), .S(n3465), .Z(N2674) );
  CMX2X1 U17586 ( .A0(mem_data1[613]), .A1(mem_data1[614]), .S(n3869), .Z(
        n8271) );
  CMXI2X1 U17587 ( .A0(n8271), .A1(n8258), .S(n4036), .Z(n8278) );
  CMX2X1 U17588 ( .A0(n8259), .A1(n8278), .S(n4351), .Z(n8291) );
  CMXI2X1 U17589 ( .A0(n8260), .A1(n8291), .S(n3465), .Z(N2675) );
  CMX2X1 U17590 ( .A0(mem_data1[73]), .A1(mem_data1[74]), .S(n3870), .Z(n8331)
         );
  CMXI2X1 U17591 ( .A0(n8331), .A1(n8261), .S(n4036), .Z(n8398) );
  CMX2X1 U17592 ( .A0(n8262), .A1(n8398), .S(n4351), .Z(n8531) );
  CMXI2X1 U17593 ( .A0(n8263), .A1(n8531), .S(n3464), .Z(N2135) );
  CMXI2X1 U17594 ( .A0(n4419), .A1(n8265), .S(n3779), .Z(n8267) );
  CMXI2X1 U17595 ( .A0(n8267), .A1(n8266), .S(n3464), .Z(N2081) );
  CMX2X1 U17596 ( .A0(mem_data1[614]), .A1(mem_data1[615]), .S(n3871), .Z(
        n8274) );
  CMXI2X1 U17597 ( .A0(n8274), .A1(n8268), .S(n4036), .Z(n8281) );
  CMX2X1 U17598 ( .A0(n8269), .A1(n8281), .S(n4351), .Z(n8294) );
  CMXI2X1 U17599 ( .A0(n8270), .A1(n8294), .S(n3464), .Z(N2676) );
  CMX2X1 U17600 ( .A0(mem_data1[615]), .A1(mem_data1[616]), .S(n3881), .Z(
        n8277) );
  CMXI2X1 U17601 ( .A0(n8277), .A1(n8271), .S(n4036), .Z(n8284) );
  CMX2X1 U17602 ( .A0(n8272), .A1(n8284), .S(n4351), .Z(n8297) );
  CMXI2X1 U17603 ( .A0(n8273), .A1(n8297), .S(n3464), .Z(N2677) );
  CMX2X1 U17604 ( .A0(mem_data1[616]), .A1(mem_data1[617]), .S(n3862), .Z(
        n8280) );
  CMXI2X1 U17605 ( .A0(n8280), .A1(n8274), .S(n4036), .Z(n8287) );
  CMX2X1 U17606 ( .A0(n8275), .A1(n8287), .S(n4351), .Z(n8303) );
  CMXI2X1 U17607 ( .A0(n8276), .A1(n8303), .S(n3467), .Z(N2678) );
  CMX2X1 U17608 ( .A0(mem_data1[617]), .A1(mem_data1[618]), .S(n3863), .Z(
        n8283) );
  CMXI2X1 U17609 ( .A0(n8283), .A1(n8277), .S(n4036), .Z(n8290) );
  CMX2X1 U17610 ( .A0(n8278), .A1(n8290), .S(n4351), .Z(n8306) );
  CMXI2X1 U17611 ( .A0(n8279), .A1(n8306), .S(n3467), .Z(N2679) );
  CMX2X1 U17612 ( .A0(mem_data1[618]), .A1(mem_data1[619]), .S(n3864), .Z(
        n8286) );
  CMXI2X1 U17613 ( .A0(n8286), .A1(n8280), .S(n4036), .Z(n8293) );
  CMX2X1 U17614 ( .A0(n8281), .A1(n8293), .S(n4351), .Z(n8309) );
  CMXI2X1 U17615 ( .A0(n8282), .A1(n8309), .S(n3467), .Z(N2680) );
  CMX2X1 U17616 ( .A0(mem_data1[619]), .A1(mem_data1[620]), .S(n3878), .Z(
        n8289) );
  CMXI2X1 U17617 ( .A0(n8289), .A1(n8283), .S(n4036), .Z(n8296) );
  CMX2X1 U17618 ( .A0(n8284), .A1(n8296), .S(n4351), .Z(n8312) );
  CMXI2X1 U17619 ( .A0(n8285), .A1(n8312), .S(n3467), .Z(N2681) );
  CMX2X1 U17620 ( .A0(mem_data1[620]), .A1(mem_data1[621]), .S(n3874), .Z(
        n8292) );
  CMXI2X1 U17621 ( .A0(n8292), .A1(n8286), .S(n4036), .Z(n8302) );
  CMX2X1 U17622 ( .A0(n8287), .A1(n8302), .S(n4351), .Z(n8315) );
  CMXI2X1 U17623 ( .A0(n8288), .A1(n8315), .S(n3467), .Z(N2682) );
  CMX2X1 U17624 ( .A0(mem_data1[621]), .A1(mem_data1[622]), .S(n3875), .Z(
        n8295) );
  CMXI2X1 U17625 ( .A0(n8295), .A1(n8289), .S(n4036), .Z(n8305) );
  CMX2X1 U17626 ( .A0(n8290), .A1(n8305), .S(n4351), .Z(n8318) );
  CMXI2X1 U17627 ( .A0(n8291), .A1(n8318), .S(n3467), .Z(N2683) );
  CMX2X1 U17628 ( .A0(mem_data1[622]), .A1(mem_data1[623]), .S(n3876), .Z(
        n8301) );
  CMXI2X1 U17629 ( .A0(n8301), .A1(n8292), .S(n4035), .Z(n8308) );
  CMX2X1 U17630 ( .A0(n8293), .A1(n8308), .S(n4351), .Z(n8321) );
  CMXI2X1 U17631 ( .A0(n8294), .A1(n8321), .S(n3467), .Z(N2684) );
  CMX2X1 U17632 ( .A0(mem_data1[623]), .A1(mem_data1[624]), .S(n3877), .Z(
        n8304) );
  CMXI2X1 U17633 ( .A0(n8304), .A1(n8295), .S(n4035), .Z(n8311) );
  CMX2X1 U17634 ( .A0(n8296), .A1(n8311), .S(n4350), .Z(n8324) );
  CMXI2X1 U17635 ( .A0(n8297), .A1(n8324), .S(n3467), .Z(N2685) );
  CMX2X1 U17636 ( .A0(mem_data1[74]), .A1(mem_data1[75]), .S(n3878), .Z(n8364)
         );
  CMXI2X1 U17637 ( .A0(n8364), .A1(n8298), .S(n4035), .Z(n8431) );
  CMX2X1 U17638 ( .A0(n8299), .A1(n8431), .S(n4350), .Z(n8564) );
  CMXI2X1 U17639 ( .A0(n8300), .A1(n8564), .S(n3467), .Z(N2136) );
  CMX2X1 U17640 ( .A0(mem_data1[624]), .A1(mem_data1[625]), .S(n3879), .Z(
        n8307) );
  CMXI2X1 U17641 ( .A0(n8307), .A1(n8301), .S(n4035), .Z(n8314) );
  CMX2X1 U17642 ( .A0(n8302), .A1(n8314), .S(n4350), .Z(n8327) );
  CMXI2X1 U17643 ( .A0(n8303), .A1(n8327), .S(n3467), .Z(N2686) );
  CMX2X1 U17644 ( .A0(mem_data1[625]), .A1(mem_data1[626]), .S(n3880), .Z(
        n8310) );
  CMXI2X1 U17645 ( .A0(n8310), .A1(n8304), .S(n4035), .Z(n8317) );
  CMX2X1 U17646 ( .A0(n8305), .A1(n8317), .S(n4350), .Z(n8330) );
  CMXI2X1 U17647 ( .A0(n8306), .A1(n8330), .S(n3466), .Z(N2687) );
  CMX2X1 U17648 ( .A0(mem_data1[626]), .A1(mem_data1[627]), .S(n3876), .Z(
        n8313) );
  CMXI2X1 U17649 ( .A0(n8313), .A1(n8307), .S(n4035), .Z(n8320) );
  CMX2X1 U17650 ( .A0(n8308), .A1(n8320), .S(n4350), .Z(n8336) );
  CMXI2X1 U17651 ( .A0(n8309), .A1(n8336), .S(n3466), .Z(N2688) );
  CMX2X1 U17652 ( .A0(mem_data1[627]), .A1(mem_data1[628]), .S(n3877), .Z(
        n8316) );
  CMXI2X1 U17653 ( .A0(n8316), .A1(n8310), .S(n4035), .Z(n8323) );
  CMX2X1 U17654 ( .A0(n8311), .A1(n8323), .S(n4350), .Z(n8339) );
  CMXI2X1 U17655 ( .A0(n8312), .A1(n8339), .S(n3466), .Z(N2689) );
  CMX2X1 U17656 ( .A0(mem_data1[628]), .A1(mem_data1[629]), .S(n3881), .Z(
        n8319) );
  CMXI2X1 U17657 ( .A0(n8319), .A1(n8313), .S(n4035), .Z(n8326) );
  CMX2X1 U17658 ( .A0(n8314), .A1(n8326), .S(n4350), .Z(n8342) );
  CMXI2X1 U17659 ( .A0(n8315), .A1(n8342), .S(n3466), .Z(N2690) );
  CMX2X1 U17660 ( .A0(mem_data1[629]), .A1(mem_data1[630]), .S(n3862), .Z(
        n8322) );
  CMXI2X1 U17661 ( .A0(n8322), .A1(n8316), .S(n4035), .Z(n8329) );
  CMX2X1 U17662 ( .A0(n8317), .A1(n8329), .S(n4350), .Z(n8345) );
  CMXI2X1 U17663 ( .A0(n8318), .A1(n8345), .S(n3466), .Z(N2691) );
  CMX2X1 U17664 ( .A0(mem_data1[630]), .A1(mem_data1[631]), .S(n3872), .Z(
        n8325) );
  CMXI2X1 U17665 ( .A0(n8325), .A1(n8319), .S(n4035), .Z(n8335) );
  CMX2X1 U17666 ( .A0(n8320), .A1(n8335), .S(n4350), .Z(n8348) );
  CMXI2X1 U17667 ( .A0(n8321), .A1(n8348), .S(n3466), .Z(N2692) );
  CMX2X1 U17668 ( .A0(mem_data1[631]), .A1(mem_data1[632]), .S(n3873), .Z(
        n8328) );
  CMXI2X1 U17669 ( .A0(n8328), .A1(n8322), .S(n4035), .Z(n8338) );
  CMX2X1 U17670 ( .A0(n8323), .A1(n8338), .S(n4350), .Z(n8351) );
  CMXI2X1 U17671 ( .A0(n8324), .A1(n8351), .S(n3466), .Z(N2693) );
  CMX2X1 U17672 ( .A0(mem_data1[632]), .A1(mem_data1[633]), .S(n3874), .Z(
        n8334) );
  CMXI2X1 U17673 ( .A0(n8334), .A1(n8325), .S(n4035), .Z(n8341) );
  CMX2X1 U17674 ( .A0(n8326), .A1(n8341), .S(n4350), .Z(n8354) );
  CMXI2X1 U17675 ( .A0(n8327), .A1(n8354), .S(n3466), .Z(N2694) );
  CMX2X1 U17676 ( .A0(mem_data1[633]), .A1(mem_data1[634]), .S(n3875), .Z(
        n8337) );
  CMXI2X1 U17677 ( .A0(n8337), .A1(n8328), .S(n4035), .Z(n8344) );
  CMX2X1 U17678 ( .A0(n8329), .A1(n8344), .S(n4349), .Z(n8357) );
  CMXI2X1 U17679 ( .A0(n8330), .A1(n8357), .S(n3469), .Z(N2695) );
  CMX2X1 U17680 ( .A0(mem_data1[75]), .A1(mem_data1[76]), .S(n3865), .Z(n8397)
         );
  CMXI2X1 U17681 ( .A0(n8397), .A1(n8331), .S(n4035), .Z(n8464) );
  CMX2X1 U17682 ( .A0(n8332), .A1(n8464), .S(n4349), .Z(n8597) );
  CMXI2X1 U17683 ( .A0(n8333), .A1(n8597), .S(n3469), .Z(N2137) );
  CMX2X1 U17684 ( .A0(mem_data1[634]), .A1(mem_data1[635]), .S(n3866), .Z(
        n8340) );
  CMXI2X1 U17685 ( .A0(n8340), .A1(n8334), .S(n4035), .Z(n8347) );
  CMX2X1 U17686 ( .A0(n8335), .A1(n8347), .S(n4349), .Z(n8360) );
  CMXI2X1 U17687 ( .A0(n8336), .A1(n8360), .S(n3469), .Z(N2696) );
  CMX2X1 U17688 ( .A0(mem_data1[635]), .A1(mem_data1[636]), .S(n3867), .Z(
        n8343) );
  CMXI2X1 U17689 ( .A0(n8343), .A1(n8337), .S(n4035), .Z(n8350) );
  CMX2X1 U17690 ( .A0(n8338), .A1(n8350), .S(n4349), .Z(n8363) );
  CMXI2X1 U17691 ( .A0(n8339), .A1(n8363), .S(n3469), .Z(N2697) );
  CMX2X1 U17692 ( .A0(mem_data1[636]), .A1(mem_data1[637]), .S(n3868), .Z(
        n8346) );
  CMXI2X1 U17693 ( .A0(n8346), .A1(n8340), .S(n4034), .Z(n8353) );
  CMX2X1 U17694 ( .A0(n8341), .A1(n8353), .S(n4349), .Z(n8369) );
  CMXI2X1 U17695 ( .A0(n8342), .A1(n8369), .S(n3469), .Z(N2698) );
  CMX2X1 U17696 ( .A0(mem_data1[637]), .A1(mem_data1[638]), .S(n3879), .Z(
        n8349) );
  CMXI2X1 U17697 ( .A0(n8349), .A1(n8343), .S(n4034), .Z(n8356) );
  CMX2X1 U17698 ( .A0(n8344), .A1(n8356), .S(n4349), .Z(n8372) );
  CMXI2X1 U17699 ( .A0(n8345), .A1(n8372), .S(n3469), .Z(N2699) );
  CMX2X1 U17700 ( .A0(mem_data1[638]), .A1(mem_data1[639]), .S(n3863), .Z(
        n8352) );
  CMXI2X1 U17701 ( .A0(n8352), .A1(n8346), .S(n4034), .Z(n8359) );
  CMX2X1 U17702 ( .A0(n8347), .A1(n8359), .S(n4349), .Z(n8375) );
  CMXI2X1 U17703 ( .A0(n8348), .A1(n8375), .S(n3468), .Z(N2700) );
  CMX2X1 U17704 ( .A0(mem_data1[639]), .A1(mem_data1[640]), .S(n3864), .Z(
        n8355) );
  CMXI2X1 U17705 ( .A0(n8355), .A1(n8349), .S(n4034), .Z(n8362) );
  CMX2X1 U17706 ( .A0(n8350), .A1(n8362), .S(n4349), .Z(n8378) );
  CMXI2X1 U17707 ( .A0(n8351), .A1(n8378), .S(n3468), .Z(N2701) );
  CMX2X1 U17708 ( .A0(mem_data1[640]), .A1(mem_data1[641]), .S(n3865), .Z(
        n8358) );
  CMXI2X1 U17709 ( .A0(n8358), .A1(n8352), .S(n4034), .Z(n8368) );
  CMX2X1 U17710 ( .A0(n8353), .A1(n8368), .S(n4349), .Z(n8381) );
  CMXI2X1 U17711 ( .A0(n8354), .A1(n8381), .S(n3468), .Z(N2702) );
  CMX2X1 U17712 ( .A0(mem_data1[641]), .A1(mem_data1[642]), .S(n3866), .Z(
        n8361) );
  CMXI2X1 U17713 ( .A0(n8361), .A1(n8355), .S(n4034), .Z(n8371) );
  CMX2X1 U17714 ( .A0(n8356), .A1(n8371), .S(n4349), .Z(n8384) );
  CMXI2X1 U17715 ( .A0(n8357), .A1(n8384), .S(n3468), .Z(N2703) );
  CMX2X1 U17716 ( .A0(mem_data1[642]), .A1(mem_data1[643]), .S(n3867), .Z(
        n8367) );
  CMXI2X1 U17717 ( .A0(n8367), .A1(n8358), .S(n4034), .Z(n8374) );
  CMX2X1 U17718 ( .A0(n8359), .A1(n8374), .S(n4349), .Z(n8387) );
  CMXI2X1 U17719 ( .A0(n8360), .A1(n8387), .S(n3468), .Z(N2704) );
  CMX2X1 U17720 ( .A0(mem_data1[643]), .A1(mem_data1[644]), .S(n3868), .Z(
        n8370) );
  CMXI2X1 U17721 ( .A0(n8370), .A1(n8361), .S(n4034), .Z(n8377) );
  CMX2X1 U17722 ( .A0(n8362), .A1(n8377), .S(n4348), .Z(n8390) );
  CMXI2X1 U17723 ( .A0(n8363), .A1(n8390), .S(n3468), .Z(N2705) );
  CMX2X1 U17724 ( .A0(mem_data1[76]), .A1(mem_data1[77]), .S(n3869), .Z(n8430)
         );
  CMXI2X1 U17725 ( .A0(n8430), .A1(n8364), .S(n4034), .Z(n8497) );
  CMX2X1 U17726 ( .A0(n8365), .A1(n8497), .S(n4348), .Z(n8634) );
  CMXI2X1 U17727 ( .A0(n8366), .A1(n8634), .S(n3468), .Z(N2138) );
  CMX2X1 U17728 ( .A0(mem_data1[644]), .A1(mem_data1[645]), .S(n3878), .Z(
        n8373) );
  CMXI2X1 U17729 ( .A0(n8373), .A1(n8367), .S(n4034), .Z(n8380) );
  CMX2X1 U17730 ( .A0(n8368), .A1(n8380), .S(n4348), .Z(n8393) );
  CMXI2X1 U17731 ( .A0(n8369), .A1(n8393), .S(n3468), .Z(N2706) );
  CMX2X1 U17732 ( .A0(mem_data1[645]), .A1(mem_data1[646]), .S(n3879), .Z(
        n8376) );
  CMXI2X1 U17733 ( .A0(n8376), .A1(n8370), .S(n4034), .Z(n8383) );
  CMX2X1 U17734 ( .A0(n8371), .A1(n8383), .S(n4348), .Z(n8396) );
  CMXI2X1 U17735 ( .A0(n8372), .A1(n8396), .S(n3468), .Z(N2707) );
  CMX2X1 U17736 ( .A0(mem_data1[646]), .A1(mem_data1[647]), .S(n3870), .Z(
        n8379) );
  CMXI2X1 U17737 ( .A0(n8379), .A1(n8373), .S(n4034), .Z(n8386) );
  CMX2X1 U17738 ( .A0(n8374), .A1(n8386), .S(n4348), .Z(n8402) );
  CMXI2X1 U17739 ( .A0(n8375), .A1(n8402), .S(n3468), .Z(N2708) );
  CMX2X1 U17740 ( .A0(mem_data1[647]), .A1(mem_data1[648]), .S(n3871), .Z(
        n8382) );
  CMXI2X1 U17741 ( .A0(n8382), .A1(n8376), .S(n4034), .Z(n8389) );
  CMX2X1 U17742 ( .A0(n8377), .A1(n8389), .S(n4348), .Z(n8405) );
  CMXI2X1 U17743 ( .A0(n8378), .A1(n8405), .S(n3468), .Z(N2709) );
  CMX2X1 U17744 ( .A0(mem_data1[648]), .A1(mem_data1[649]), .S(n3876), .Z(
        n8385) );
  CMXI2X1 U17745 ( .A0(n8385), .A1(n8379), .S(n4034), .Z(n8392) );
  CMX2X1 U17746 ( .A0(n8380), .A1(n8392), .S(n4348), .Z(n8408) );
  CMXI2X1 U17747 ( .A0(n8381), .A1(n8408), .S(n3467), .Z(N2710) );
  CMX2X1 U17748 ( .A0(mem_data1[649]), .A1(mem_data1[650]), .S(n3877), .Z(
        n8388) );
  CMXI2X1 U17749 ( .A0(n8388), .A1(n8382), .S(n4034), .Z(n8395) );
  CMX2X1 U17750 ( .A0(n8383), .A1(n8395), .S(n4348), .Z(n8411) );
  CMXI2X1 U17751 ( .A0(n8384), .A1(n8411), .S(n3471), .Z(N2711) );
  CMX2X1 U17752 ( .A0(mem_data1[650]), .A1(mem_data1[651]), .S(n3878), .Z(
        n8391) );
  CMXI2X1 U17753 ( .A0(n8391), .A1(n8385), .S(n4034), .Z(n8401) );
  CMX2X1 U17754 ( .A0(n8386), .A1(n8401), .S(n4348), .Z(n8414) );
  CMXI2X1 U17755 ( .A0(n8387), .A1(n8414), .S(n3471), .Z(N2712) );
  CMX2X1 U17756 ( .A0(mem_data1[651]), .A1(mem_data1[652]), .S(n3879), .Z(
        n8394) );
  CMXI2X1 U17757 ( .A0(n8394), .A1(n8388), .S(n4033), .Z(n8404) );
  CMX2X1 U17758 ( .A0(n8389), .A1(n8404), .S(n4348), .Z(n8417) );
  CMXI2X1 U17759 ( .A0(n8390), .A1(n8417), .S(n3470), .Z(N2713) );
  CMX2X1 U17760 ( .A0(mem_data1[652]), .A1(mem_data1[653]), .S(n3869), .Z(
        n8400) );
  CMXI2X1 U17761 ( .A0(n8400), .A1(n8391), .S(n4033), .Z(n8407) );
  CMX2X1 U17762 ( .A0(n8392), .A1(n8407), .S(n4348), .Z(n8420) );
  CMXI2X1 U17763 ( .A0(n8393), .A1(n8420), .S(n3470), .Z(N2714) );
  CMX2X1 U17764 ( .A0(mem_data1[653]), .A1(mem_data1[654]), .S(n3870), .Z(
        n8403) );
  CMXI2X1 U17765 ( .A0(n8403), .A1(n8394), .S(n4033), .Z(n8410) );
  CMX2X1 U17766 ( .A0(n8395), .A1(n8410), .S(n4347), .Z(n8423) );
  CMXI2X1 U17767 ( .A0(n8396), .A1(n8423), .S(n3470), .Z(N2715) );
  CMX2X1 U17768 ( .A0(mem_data1[77]), .A1(mem_data1[78]), .S(n3871), .Z(n8463)
         );
  CMXI2X1 U17769 ( .A0(n8463), .A1(n8397), .S(n4033), .Z(n8530) );
  CMX2X1 U17770 ( .A0(n8398), .A1(n8530), .S(n4347), .Z(n8667) );
  CMXI2X1 U17771 ( .A0(n8399), .A1(n8667), .S(n3470), .Z(N2139) );
  CMX2X1 U17772 ( .A0(mem_data1[654]), .A1(mem_data1[655]), .S(n3872), .Z(
        n8406) );
  CMXI2X1 U17773 ( .A0(n8406), .A1(n8400), .S(n4033), .Z(n8413) );
  CMX2X1 U17774 ( .A0(n8401), .A1(n8413), .S(n4347), .Z(n8426) );
  CMXI2X1 U17775 ( .A0(n8402), .A1(n8426), .S(n3470), .Z(N2716) );
  CMX2X1 U17776 ( .A0(mem_data1[655]), .A1(mem_data1[656]), .S(n3880), .Z(
        n8409) );
  CMXI2X1 U17777 ( .A0(n8409), .A1(n8403), .S(n4033), .Z(n8416) );
  CMX2X1 U17778 ( .A0(n8404), .A1(n8416), .S(n4347), .Z(n8429) );
  CMXI2X1 U17779 ( .A0(n8405), .A1(n8429), .S(n3470), .Z(N2717) );
  CMX2X1 U17780 ( .A0(mem_data1[656]), .A1(mem_data1[657]), .S(n3872), .Z(
        n8412) );
  CMXI2X1 U17781 ( .A0(n8412), .A1(n8406), .S(n4033), .Z(n8419) );
  CMX2X1 U17782 ( .A0(n8407), .A1(n8419), .S(n4347), .Z(n8435) );
  CMXI2X1 U17783 ( .A0(n8408), .A1(n8435), .S(n3470), .Z(N2718) );
  CMX2X1 U17784 ( .A0(mem_data1[657]), .A1(mem_data1[658]), .S(n3873), .Z(
        n8415) );
  CMXI2X1 U17785 ( .A0(n8415), .A1(n8409), .S(n4033), .Z(n8422) );
  CMX2X1 U17786 ( .A0(n8410), .A1(n8422), .S(n4347), .Z(n8438) );
  CMXI2X1 U17787 ( .A0(n8411), .A1(n8438), .S(n3470), .Z(N2719) );
  CMX2X1 U17788 ( .A0(mem_data1[658]), .A1(mem_data1[659]), .S(n3874), .Z(
        n8418) );
  CMXI2X1 U17789 ( .A0(n8418), .A1(n8412), .S(n4033), .Z(n8425) );
  CMX2X1 U17790 ( .A0(n8413), .A1(n8425), .S(n4347), .Z(n8441) );
  CMXI2X1 U17791 ( .A0(n8414), .A1(n8441), .S(n3470), .Z(N2720) );
  CMX2X1 U17792 ( .A0(mem_data1[659]), .A1(mem_data1[660]), .S(n3875), .Z(
        n8421) );
  CMXI2X1 U17793 ( .A0(n8421), .A1(n8415), .S(n4033), .Z(n8428) );
  CMX2X1 U17794 ( .A0(n8416), .A1(n8428), .S(n4347), .Z(n8444) );
  CMXI2X1 U17795 ( .A0(n8417), .A1(n8444), .S(n3470), .Z(N2721) );
  CMX2X1 U17796 ( .A0(mem_data1[660]), .A1(mem_data1[661]), .S(n3876), .Z(
        n8424) );
  CMXI2X1 U17797 ( .A0(n8424), .A1(n8418), .S(n4033), .Z(n8434) );
  CMX2X1 U17798 ( .A0(n8419), .A1(n8434), .S(n4347), .Z(n8447) );
  CMXI2X1 U17799 ( .A0(n8420), .A1(n8447), .S(n3470), .Z(N2722) );
  CMX2X1 U17800 ( .A0(mem_data1[661]), .A1(mem_data1[662]), .S(n3877), .Z(
        n8427) );
  CMXI2X1 U17801 ( .A0(n8427), .A1(n8421), .S(n4033), .Z(n8437) );
  CMX2X1 U17802 ( .A0(n8422), .A1(n8437), .S(n4347), .Z(n8450) );
  CMXI2X1 U17803 ( .A0(n8423), .A1(n8450), .S(n3469), .Z(N2723) );
  CMX2X1 U17804 ( .A0(mem_data1[662]), .A1(mem_data1[663]), .S(n3878), .Z(
        n8433) );
  CMXI2X1 U17805 ( .A0(n8433), .A1(n8424), .S(n4033), .Z(n8440) );
  CMX2X1 U17806 ( .A0(n8425), .A1(n8440), .S(n4347), .Z(n8453) );
  CMXI2X1 U17807 ( .A0(n8426), .A1(n8453), .S(n3469), .Z(N2724) );
  CMX2X1 U17808 ( .A0(mem_data1[663]), .A1(mem_data1[664]), .S(n3880), .Z(
        n8436) );
  CMXI2X1 U17809 ( .A0(n8436), .A1(n8427), .S(n4033), .Z(n8443) );
  CMX2X1 U17810 ( .A0(n8428), .A1(n8443), .S(n4346), .Z(n8456) );
  CMXI2X1 U17811 ( .A0(n8429), .A1(n8456), .S(n3469), .Z(N2725) );
  CMX2X1 U17812 ( .A0(mem_data1[78]), .A1(mem_data1[79]), .S(n3881), .Z(n8496)
         );
  CMXI2X1 U17813 ( .A0(n8496), .A1(n8430), .S(n4033), .Z(n8563) );
  CMX2X1 U17814 ( .A0(n8431), .A1(n8563), .S(n4346), .Z(n8700) );
  CMXI2X1 U17815 ( .A0(n8432), .A1(n8700), .S(n3469), .Z(N2140) );
  CMX2X1 U17816 ( .A0(mem_data1[664]), .A1(mem_data1[665]), .S(n3879), .Z(
        n8439) );
  CMXI2X1 U17817 ( .A0(n8439), .A1(n8433), .S(n4033), .Z(n8446) );
  CMX2X1 U17818 ( .A0(n8434), .A1(n8446), .S(n4346), .Z(n8459) );
  CMXI2X1 U17819 ( .A0(n8435), .A1(n8459), .S(n3469), .Z(N2726) );
  CMX2X1 U17820 ( .A0(mem_data1[665]), .A1(mem_data1[666]), .S(n3880), .Z(
        n8442) );
  CMXI2X1 U17821 ( .A0(n8442), .A1(n8436), .S(n4032), .Z(n8449) );
  CMX2X1 U17822 ( .A0(n8437), .A1(n8449), .S(n4346), .Z(n8462) );
  CMXI2X1 U17823 ( .A0(n8438), .A1(n8462), .S(n3472), .Z(N2727) );
  CMX2X1 U17824 ( .A0(mem_data1[666]), .A1(mem_data1[667]), .S(n3880), .Z(
        n8445) );
  CMXI2X1 U17825 ( .A0(n8445), .A1(n8439), .S(n4032), .Z(n8452) );
  CMX2X1 U17826 ( .A0(n8440), .A1(n8452), .S(n4346), .Z(n8468) );
  CMXI2X1 U17827 ( .A0(n8441), .A1(n8468), .S(n3472), .Z(N2728) );
  CMX2X1 U17828 ( .A0(mem_data1[667]), .A1(mem_data1[668]), .S(n3881), .Z(
        n8448) );
  CMXI2X1 U17829 ( .A0(n8448), .A1(n8442), .S(n4032), .Z(n8455) );
  CMX2X1 U17830 ( .A0(n8443), .A1(n8455), .S(n4346), .Z(n8471) );
  CMXI2X1 U17831 ( .A0(n8444), .A1(n8471), .S(n3472), .Z(N2729) );
  CMX2X1 U17832 ( .A0(mem_data1[668]), .A1(mem_data1[669]), .S(n3862), .Z(
        n8451) );
  CMXI2X1 U17833 ( .A0(n8451), .A1(n8445), .S(n4032), .Z(n8458) );
  CMX2X1 U17834 ( .A0(n8446), .A1(n8458), .S(n4346), .Z(n8474) );
  CMXI2X1 U17835 ( .A0(n8447), .A1(n8474), .S(n3472), .Z(N2730) );
  CMX2X1 U17836 ( .A0(mem_data1[669]), .A1(mem_data1[670]), .S(n3863), .Z(
        n8454) );
  CMXI2X1 U17837 ( .A0(n8454), .A1(n8448), .S(n4032), .Z(n8461) );
  CMX2X1 U17838 ( .A0(n8449), .A1(n8461), .S(n4346), .Z(n8477) );
  CMXI2X1 U17839 ( .A0(n8450), .A1(n8477), .S(n3472), .Z(N2731) );
  CMX2X1 U17840 ( .A0(mem_data1[670]), .A1(mem_data1[671]), .S(n3873), .Z(
        n8457) );
  CMXI2X1 U17841 ( .A0(n8457), .A1(n8451), .S(n4032), .Z(n8467) );
  CMX2X1 U17842 ( .A0(n8452), .A1(n8467), .S(n4346), .Z(n8480) );
  CMXI2X1 U17843 ( .A0(n8453), .A1(n8480), .S(n3472), .Z(N2732) );
  CMX2X1 U17844 ( .A0(mem_data1[671]), .A1(mem_data1[672]), .S(n3874), .Z(
        n8460) );
  CMXI2X1 U17845 ( .A0(n8460), .A1(n8454), .S(n4032), .Z(n8470) );
  CMX2X1 U17846 ( .A0(n8455), .A1(n8470), .S(n4346), .Z(n8483) );
  CMXI2X1 U17847 ( .A0(n8456), .A1(n8483), .S(n3472), .Z(N2733) );
  CMX2X1 U17848 ( .A0(mem_data1[672]), .A1(mem_data1[673]), .S(n3876), .Z(
        n8466) );
  CMXI2X1 U17849 ( .A0(n8466), .A1(n8457), .S(n4032), .Z(n8473) );
  CMX2X1 U17850 ( .A0(n8458), .A1(n8473), .S(n4346), .Z(n8486) );
  CMXI2X1 U17851 ( .A0(n8459), .A1(n8486), .S(n3472), .Z(N2734) );
  CMX2X1 U17852 ( .A0(mem_data1[673]), .A1(mem_data1[674]), .S(n3881), .Z(
        n8469) );
  CMXI2X1 U17853 ( .A0(n8469), .A1(n8460), .S(n4032), .Z(n8476) );
  CMX2X1 U17854 ( .A0(n8461), .A1(n8476), .S(n4345), .Z(n8489) );
  CMXI2X1 U17855 ( .A0(n8462), .A1(n8489), .S(n3472), .Z(N2735) );
  CMX2X1 U17856 ( .A0(mem_data1[79]), .A1(mem_data1[80]), .S(n3881), .Z(n8529)
         );
  CMXI2X1 U17857 ( .A0(n8529), .A1(n8463), .S(n4032), .Z(n8596) );
  CMX2X1 U17858 ( .A0(n8464), .A1(n8596), .S(n4345), .Z(n8733) );
  CMXI2X1 U17859 ( .A0(n8465), .A1(n8733), .S(n3471), .Z(N2141) );
  CMX2X1 U17860 ( .A0(mem_data1[674]), .A1(mem_data1[675]), .S(n3862), .Z(
        n8472) );
  CMXI2X1 U17861 ( .A0(n8472), .A1(n8466), .S(n4032), .Z(n8479) );
  CMX2X1 U17862 ( .A0(n8467), .A1(n8479), .S(n4345), .Z(n8492) );
  CMXI2X1 U17863 ( .A0(n8468), .A1(n8492), .S(n3471), .Z(N2736) );
  CMX2X1 U17864 ( .A0(mem_data1[675]), .A1(mem_data1[676]), .S(n3863), .Z(
        n8475) );
  CMXI2X1 U17865 ( .A0(n8475), .A1(n8469), .S(n4032), .Z(n8482) );
  CMX2X1 U17866 ( .A0(n8470), .A1(n8482), .S(n4345), .Z(n8495) );
  CMXI2X1 U17867 ( .A0(n8471), .A1(n8495), .S(n3471), .Z(N2737) );
  CMX2X1 U17868 ( .A0(mem_data1[676]), .A1(mem_data1[677]), .S(n3864), .Z(
        n8478) );
  CMXI2X1 U17869 ( .A0(n8478), .A1(n8472), .S(n4032), .Z(n8485) );
  CMX2X1 U17870 ( .A0(n8473), .A1(n8485), .S(n4345), .Z(n8501) );
  CMXI2X1 U17871 ( .A0(n8474), .A1(n8501), .S(n3471), .Z(N2738) );
  CMX2X1 U17872 ( .A0(mem_data1[677]), .A1(mem_data1[678]), .S(n3865), .Z(
        n8481) );
  CMXI2X1 U17873 ( .A0(n8481), .A1(n8475), .S(n4032), .Z(n8488) );
  CMX2X1 U17874 ( .A0(n8476), .A1(n8488), .S(n4345), .Z(n8504) );
  CMXI2X1 U17875 ( .A0(n8477), .A1(n8504), .S(n3471), .Z(N2739) );
  CMX2X1 U17876 ( .A0(mem_data1[678]), .A1(mem_data1[679]), .S(n3866), .Z(
        n8484) );
  CMXI2X1 U17877 ( .A0(n8484), .A1(n8478), .S(n4032), .Z(n8491) );
  CMX2X1 U17878 ( .A0(n8479), .A1(n8491), .S(n4345), .Z(n8507) );
  CMXI2X1 U17879 ( .A0(n8480), .A1(n8507), .S(n3471), .Z(N2740) );
  CMX2X1 U17880 ( .A0(mem_data1[679]), .A1(mem_data1[680]), .S(n3867), .Z(
        n8487) );
  CMXI2X1 U17881 ( .A0(n8487), .A1(n8481), .S(n4032), .Z(n8494) );
  CMX2X1 U17882 ( .A0(n8482), .A1(n8494), .S(n4345), .Z(n8510) );
  CMXI2X1 U17883 ( .A0(n8483), .A1(n8510), .S(n3471), .Z(N2741) );
  CMX2X1 U17884 ( .A0(mem_data1[680]), .A1(mem_data1[681]), .S(n3862), .Z(
        n8490) );
  CMXI2X1 U17885 ( .A0(n8490), .A1(n8484), .S(n4031), .Z(n8500) );
  CMX2X1 U17886 ( .A0(n8485), .A1(n8500), .S(n4345), .Z(n8513) );
  CMXI2X1 U17887 ( .A0(n8486), .A1(n8513), .S(n3471), .Z(N2742) );
  CMX2X1 U17888 ( .A0(mem_data1[681]), .A1(mem_data1[682]), .S(n3863), .Z(
        n8493) );
  CMXI2X1 U17889 ( .A0(n8493), .A1(n8487), .S(n4031), .Z(n8503) );
  CMX2X1 U17890 ( .A0(n8488), .A1(n8503), .S(n4345), .Z(n8516) );
  CMXI2X1 U17891 ( .A0(n8489), .A1(n8516), .S(n3471), .Z(N2743) );
  CMX2X1 U17892 ( .A0(mem_data1[682]), .A1(mem_data1[683]), .S(n3868), .Z(
        n8499) );
  CMXI2X1 U17893 ( .A0(n8499), .A1(n8490), .S(n4031), .Z(n8506) );
  CMX2X1 U17894 ( .A0(n8491), .A1(n8506), .S(n4345), .Z(n8519) );
  CMXI2X1 U17895 ( .A0(n8492), .A1(n8519), .S(n3474), .Z(N2744) );
  CMX2X1 U17896 ( .A0(mem_data1[683]), .A1(mem_data1[684]), .S(n3869), .Z(
        n8502) );
  CMXI2X1 U17897 ( .A0(n8502), .A1(n8493), .S(n4031), .Z(n8509) );
  CMX2X1 U17898 ( .A0(n8494), .A1(n8509), .S(n4344), .Z(n8522) );
  CMXI2X1 U17899 ( .A0(n8495), .A1(n8522), .S(n3474), .Z(N2745) );
  CMX2X1 U17900 ( .A0(mem_data1[80]), .A1(mem_data1[81]), .S(n3864), .Z(n8562)
         );
  CMXI2X1 U17901 ( .A0(n8562), .A1(n8496), .S(n4031), .Z(n8633) );
  CMX2X1 U17902 ( .A0(n8497), .A1(n8633), .S(n4346), .Z(n8766) );
  CMXI2X1 U17903 ( .A0(n8498), .A1(n8766), .S(n3474), .Z(N2142) );
  CMX2X1 U17904 ( .A0(mem_data1[684]), .A1(mem_data1[685]), .S(n3865), .Z(
        n8505) );
  CMXI2X1 U17905 ( .A0(n8505), .A1(n8499), .S(n4031), .Z(n8512) );
  CMX2X1 U17906 ( .A0(n8500), .A1(n8512), .S(n4347), .Z(n8525) );
  CMXI2X1 U17907 ( .A0(n8501), .A1(n8525), .S(n3474), .Z(N2746) );
  CMX2X1 U17908 ( .A0(mem_data1[685]), .A1(mem_data1[686]), .S(n3866), .Z(
        n8508) );
  CMXI2X1 U17909 ( .A0(n8508), .A1(n8502), .S(n4031), .Z(n8515) );
  CMX2X1 U17910 ( .A0(n8503), .A1(n8515), .S(n4348), .Z(n8528) );
  CMXI2X1 U17911 ( .A0(n8504), .A1(n8528), .S(n3474), .Z(N2747) );
  CMX2X1 U17912 ( .A0(mem_data1[686]), .A1(mem_data1[687]), .S(n3867), .Z(
        n8511) );
  CMXI2X1 U17913 ( .A0(n8511), .A1(n8505), .S(n4031), .Z(n8518) );
  CMX2X1 U17914 ( .A0(n8506), .A1(n8518), .S(n4343), .Z(n8534) );
  CMXI2X1 U17915 ( .A0(n8507), .A1(n8534), .S(n3474), .Z(N2748) );
  CMX2X1 U17916 ( .A0(mem_data1[687]), .A1(mem_data1[688]), .S(n3877), .Z(
        n8514) );
  CMXI2X1 U17917 ( .A0(n8514), .A1(n8508), .S(n4031), .Z(n8521) );
  CMX2X1 U17918 ( .A0(n8509), .A1(n8521), .S(n4349), .Z(n8537) );
  CMXI2X1 U17919 ( .A0(n8510), .A1(n8537), .S(n3473), .Z(N2749) );
  CMX2X1 U17920 ( .A0(mem_data1[688]), .A1(mem_data1[689]), .S(n3878), .Z(
        n8517) );
  CMXI2X1 U17921 ( .A0(n8517), .A1(n8511), .S(n4031), .Z(n8524) );
  CMX2X1 U17922 ( .A0(n8512), .A1(n8524), .S(n4350), .Z(n8540) );
  CMXI2X1 U17923 ( .A0(n8513), .A1(n8540), .S(n3473), .Z(N2750) );
  CMX2X1 U17924 ( .A0(mem_data1[689]), .A1(mem_data1[690]), .S(n3879), .Z(
        n8520) );
  CMXI2X1 U17925 ( .A0(n8520), .A1(n8514), .S(n4031), .Z(n8527) );
  CMX2X1 U17926 ( .A0(n8515), .A1(n8527), .S(n4351), .Z(n8543) );
  CMXI2X1 U17927 ( .A0(n8516), .A1(n8543), .S(n3473), .Z(N2751) );
  CMX2X1 U17928 ( .A0(mem_data1[690]), .A1(mem_data1[691]), .S(n3880), .Z(
        n8523) );
  CMXI2X1 U17929 ( .A0(n8523), .A1(n8517), .S(n4031), .Z(n8533) );
  CMX2X1 U17930 ( .A0(n8518), .A1(n8533), .S(n4345), .Z(n8546) );
  CMXI2X1 U17931 ( .A0(n8519), .A1(n8546), .S(n3473), .Z(N2752) );
  CMX2X1 U17932 ( .A0(mem_data1[691]), .A1(mem_data1[692]), .S(n3862), .Z(
        n8526) );
  CMXI2X1 U17933 ( .A0(n8526), .A1(n8520), .S(n4031), .Z(n8536) );
  CMX2X1 U17934 ( .A0(n8521), .A1(n8536), .S(n4341), .Z(n8549) );
  CMXI2X1 U17935 ( .A0(n8522), .A1(n8549), .S(n3473), .Z(N2753) );
  CMX2X1 U17936 ( .A0(mem_data1[692]), .A1(mem_data1[693]), .S(n3870), .Z(
        n8532) );
  CMXI2X1 U17937 ( .A0(n8532), .A1(n8523), .S(n4031), .Z(n8539) );
  CMX2X1 U17938 ( .A0(n8524), .A1(n8539), .S(n4344), .Z(n8552) );
  CMXI2X1 U17939 ( .A0(n8525), .A1(n8552), .S(n3473), .Z(N2754) );
  CMX2X1 U17940 ( .A0(mem_data1[693]), .A1(mem_data1[694]), .S(n3871), .Z(
        n8535) );
  CMXI2X1 U17941 ( .A0(n8535), .A1(n8526), .S(n4031), .Z(n8542) );
  CMX2X1 U17942 ( .A0(n8527), .A1(n8542), .S(n4344), .Z(n8555) );
  CMXI2X1 U17943 ( .A0(n8528), .A1(n8555), .S(n3473), .Z(N2755) );
  CMX2X1 U17944 ( .A0(mem_data1[81]), .A1(mem_data1[82]), .S(n3872), .Z(n8595)
         );
  CMXI2X1 U17945 ( .A0(n8595), .A1(n8529), .S(n4031), .Z(n8666) );
  CMX2X1 U17946 ( .A0(n8530), .A1(n8666), .S(n4344), .Z(n8799) );
  CMXI2X1 U17947 ( .A0(n8531), .A1(n8799), .S(n3473), .Z(N2143) );
  CMX2X1 U17948 ( .A0(mem_data1[694]), .A1(mem_data1[695]), .S(n3873), .Z(
        n8538) );
  CMXI2X1 U17949 ( .A0(n8538), .A1(n8532), .S(n4030), .Z(n8545) );
  CMX2X1 U17950 ( .A0(n8533), .A1(n8545), .S(n4344), .Z(n8558) );
  CMXI2X1 U17951 ( .A0(n8534), .A1(n8558), .S(n3473), .Z(N2756) );
  CMX2X1 U17952 ( .A0(mem_data1[695]), .A1(mem_data1[696]), .S(n3874), .Z(
        n8541) );
  CMXI2X1 U17953 ( .A0(n8541), .A1(n8535), .S(n4030), .Z(n8548) );
  CMX2X1 U17954 ( .A0(n8536), .A1(n8548), .S(n4344), .Z(n8561) );
  CMXI2X1 U17955 ( .A0(n8537), .A1(n8561), .S(n3473), .Z(N2757) );
  CMX2X1 U17956 ( .A0(mem_data1[696]), .A1(mem_data1[697]), .S(n3875), .Z(
        n8544) );
  CMXI2X1 U17957 ( .A0(n8544), .A1(n8538), .S(n4030), .Z(n8551) );
  CMX2X1 U17958 ( .A0(n8539), .A1(n8551), .S(n4344), .Z(n8567) );
  CMXI2X1 U17959 ( .A0(n8540), .A1(n8567), .S(n3472), .Z(N2758) );
  CMX2X1 U17960 ( .A0(mem_data1[697]), .A1(mem_data1[698]), .S(n3876), .Z(
        n8547) );
  CMXI2X1 U17961 ( .A0(n8547), .A1(n8541), .S(n4030), .Z(n8554) );
  CMX2X1 U17962 ( .A0(n8542), .A1(n8554), .S(n4344), .Z(n8570) );
  CMXI2X1 U17963 ( .A0(n8543), .A1(n8570), .S(n3476), .Z(N2759) );
  CMX2X1 U17964 ( .A0(mem_data1[698]), .A1(mem_data1[699]), .S(n3864), .Z(
        n8550) );
  CMXI2X1 U17965 ( .A0(n8550), .A1(n8544), .S(n4030), .Z(n8557) );
  CMX2X1 U17966 ( .A0(n8545), .A1(n8557), .S(n4344), .Z(n8573) );
  CMXI2X1 U17967 ( .A0(n8546), .A1(n8573), .S(n3476), .Z(N2760) );
  CMX2X1 U17968 ( .A0(mem_data1[699]), .A1(mem_data1[700]), .S(n3865), .Z(
        n8553) );
  CMXI2X1 U17969 ( .A0(n8553), .A1(n8547), .S(n4030), .Z(n8560) );
  CMX2X1 U17970 ( .A0(n8548), .A1(n8560), .S(n4344), .Z(n8576) );
  CMXI2X1 U17971 ( .A0(n8549), .A1(n8576), .S(n3475), .Z(N2761) );
  CMX2X1 U17972 ( .A0(mem_data1[700]), .A1(mem_data1[701]), .S(n3877), .Z(
        n8556) );
  CMXI2X1 U17973 ( .A0(n8556), .A1(n8550), .S(n4030), .Z(n8566) );
  CMX2X1 U17974 ( .A0(n8551), .A1(n8566), .S(n4344), .Z(n8579) );
  CMXI2X1 U17975 ( .A0(n8552), .A1(n8579), .S(n3475), .Z(N2762) );
  CMX2X1 U17976 ( .A0(mem_data1[701]), .A1(mem_data1[702]), .S(n3878), .Z(
        n8559) );
  CMXI2X1 U17977 ( .A0(n8559), .A1(n8553), .S(n4030), .Z(n8569) );
  CMX2X1 U17978 ( .A0(n8554), .A1(n8569), .S(n4344), .Z(n8582) );
  CMXI2X1 U17979 ( .A0(n8555), .A1(n8582), .S(n3475), .Z(N2763) );
  CMX2X1 U17980 ( .A0(mem_data1[702]), .A1(mem_data1[703]), .S(n3868), .Z(
        n8565) );
  CMXI2X1 U17981 ( .A0(n8565), .A1(n8556), .S(n4030), .Z(n8572) );
  CMX2X1 U17982 ( .A0(n8557), .A1(n8572), .S(n4343), .Z(n8585) );
  CMXI2X1 U17983 ( .A0(n8558), .A1(n8585), .S(n3475), .Z(N2764) );
  CMX2X1 U17984 ( .A0(mem_data1[703]), .A1(mem_data1[704]), .S(n3869), .Z(
        n8568) );
  CMXI2X1 U17985 ( .A0(n8568), .A1(n8559), .S(n4030), .Z(n8575) );
  CMX2X1 U17986 ( .A0(n8560), .A1(n8575), .S(n4343), .Z(n8588) );
  CMXI2X1 U17987 ( .A0(n8561), .A1(n8588), .S(n3475), .Z(N2765) );
  CMX2X1 U17988 ( .A0(mem_data1[82]), .A1(mem_data1[83]), .S(n3870), .Z(n8632)
         );
  CMXI2X1 U17989 ( .A0(n8632), .A1(n8562), .S(n4030), .Z(n8699) );
  CMX2X1 U17990 ( .A0(n8563), .A1(n8699), .S(n4343), .Z(n8832) );
  CMXI2X1 U17991 ( .A0(n8564), .A1(n8832), .S(n3475), .Z(N2144) );
  CMX2X1 U17992 ( .A0(mem_data1[704]), .A1(mem_data1[705]), .S(n3871), .Z(
        n8571) );
  CMXI2X1 U17993 ( .A0(n8571), .A1(n8565), .S(n4030), .Z(n8578) );
  CMX2X1 U17994 ( .A0(n8566), .A1(n8578), .S(n4343), .Z(n8591) );
  CMXI2X1 U17995 ( .A0(n8567), .A1(n8591), .S(n3475), .Z(N2766) );
  CMX2X1 U17996 ( .A0(mem_data1[705]), .A1(mem_data1[706]), .S(n3881), .Z(
        n8574) );
  CMXI2X1 U17997 ( .A0(n8574), .A1(n8568), .S(n4030), .Z(n8581) );
  CMX2X1 U17998 ( .A0(n8569), .A1(n8581), .S(n4343), .Z(n8594) );
  CMXI2X1 U17999 ( .A0(n8570), .A1(n8594), .S(n3475), .Z(N2767) );
  CMX2X1 U18000 ( .A0(mem_data1[706]), .A1(mem_data1[707]), .S(n3862), .Z(
        n8577) );
  CMXI2X1 U18001 ( .A0(n8577), .A1(n8571), .S(n4030), .Z(n8584) );
  CMX2X1 U18002 ( .A0(n8572), .A1(n8584), .S(n4343), .Z(n8604) );
  CMXI2X1 U18003 ( .A0(n8573), .A1(n8604), .S(n3475), .Z(N2768) );
  CMX2X1 U18004 ( .A0(mem_data1[707]), .A1(mem_data1[708]), .S(n3863), .Z(
        n8580) );
  CMXI2X1 U18005 ( .A0(n8580), .A1(n8574), .S(n4030), .Z(n8587) );
  CMX2X1 U18006 ( .A0(n8575), .A1(n8587), .S(n4343), .Z(n8607) );
  CMXI2X1 U18007 ( .A0(n8576), .A1(n8607), .S(n3475), .Z(N2769) );
  CMX2X1 U18008 ( .A0(mem_data1[708]), .A1(mem_data1[709]), .S(n3864), .Z(
        n8583) );
  CMXI2X1 U18009 ( .A0(n8583), .A1(n8577), .S(n4030), .Z(n8590) );
  CMX2X1 U18010 ( .A0(n8578), .A1(n8590), .S(n4343), .Z(n8610) );
  CMXI2X1 U18011 ( .A0(n8579), .A1(n8610), .S(n3475), .Z(N2770) );
  CMX2X1 U18012 ( .A0(mem_data1[709]), .A1(mem_data1[710]), .S(n3863), .Z(
        n8586) );
  CMXI2X1 U18013 ( .A0(n8586), .A1(n8580), .S(n4029), .Z(n8593) );
  CMX2X1 U18014 ( .A0(n8581), .A1(n8593), .S(n4343), .Z(n8613) );
  CMXI2X1 U18015 ( .A0(n8582), .A1(n8613), .S(n3474), .Z(N2771) );
  CMX2X1 U18016 ( .A0(mem_data1[710]), .A1(mem_data1[711]), .S(n3879), .Z(
        n8589) );
  CMXI2X1 U18017 ( .A0(n8589), .A1(n8583), .S(n4029), .Z(n8603) );
  CMX2X1 U18018 ( .A0(n8584), .A1(n8603), .S(n4343), .Z(n8616) );
  CMXI2X1 U18019 ( .A0(n8585), .A1(n8616), .S(n3474), .Z(N2772) );
  CMX2X1 U18020 ( .A0(mem_data1[711]), .A1(mem_data1[712]), .S(n3880), .Z(
        n8592) );
  CMXI2X1 U18021 ( .A0(n8592), .A1(n8586), .S(n4029), .Z(n8606) );
  CMX2X1 U18022 ( .A0(n8587), .A1(n8606), .S(n4343), .Z(n8619) );
  CMXI2X1 U18023 ( .A0(n8588), .A1(n8619), .S(n3474), .Z(N2773) );
  CMX2X1 U18024 ( .A0(mem_data1[712]), .A1(mem_data1[713]), .S(n3881), .Z(
        n8602) );
  CMXI2X1 U18025 ( .A0(n8602), .A1(n8589), .S(n4029), .Z(n8609) );
  CMX2X1 U18026 ( .A0(n8590), .A1(n8609), .S(n4342), .Z(n8622) );
  CMXI2X1 U18027 ( .A0(n8591), .A1(n8622), .S(n3474), .Z(N2774) );
  CMX2X1 U18028 ( .A0(mem_data1[713]), .A1(mem_data1[714]), .S(n3862), .Z(
        n8605) );
  CMXI2X1 U18029 ( .A0(n8605), .A1(n8592), .S(n4029), .Z(n8612) );
  CMX2X1 U18030 ( .A0(n8593), .A1(n8612), .S(n4342), .Z(n8625) );
  CMXI2X1 U18031 ( .A0(n8594), .A1(n8625), .S(n3474), .Z(N2775) );
  CMX2X1 U18032 ( .A0(mem_data1[83]), .A1(mem_data1[84]), .S(n3863), .Z(n8665)
         );
  CMXI2X1 U18033 ( .A0(n8665), .A1(n8595), .S(n4029), .Z(n8732) );
  CMX2X1 U18034 ( .A0(n8596), .A1(n8732), .S(n4342), .Z(n8865) );
  CMXI2X1 U18035 ( .A0(n8597), .A1(n8865), .S(n3477), .Z(N2145) );
  CMXI2X1 U18036 ( .A0(n4417), .A1(n8599), .S(n3778), .Z(n8601) );
  CMXI2X1 U18037 ( .A0(n8601), .A1(n8600), .S(n3477), .Z(N2082) );
  CMX2X1 U18038 ( .A0(mem_data1[714]), .A1(mem_data1[715]), .S(n3864), .Z(
        n8608) );
  CMXI2X1 U18039 ( .A0(n8608), .A1(n8602), .S(n4029), .Z(n8615) );
  CMX2X1 U18040 ( .A0(n8603), .A1(n8615), .S(n4342), .Z(n8628) );
  CMXI2X1 U18041 ( .A0(n8604), .A1(n8628), .S(n3477), .Z(N2776) );
  CMX2X1 U18042 ( .A0(mem_data1[715]), .A1(mem_data1[716]), .S(n3865), .Z(
        n8611) );
  CMXI2X1 U18043 ( .A0(n8611), .A1(n8605), .S(n4029), .Z(n8618) );
  CMX2X1 U18044 ( .A0(n8606), .A1(n8618), .S(n4342), .Z(n8631) );
  CMXI2X1 U18045 ( .A0(n8607), .A1(n8631), .S(n3477), .Z(N2777) );
  CMX2X1 U18046 ( .A0(mem_data1[716]), .A1(mem_data1[717]), .S(n3866), .Z(
        n8614) );
  CMXI2X1 U18047 ( .A0(n8614), .A1(n8608), .S(n4029), .Z(n8621) );
  CMX2X1 U18048 ( .A0(n8609), .A1(n8621), .S(n4342), .Z(n8637) );
  CMXI2X1 U18049 ( .A0(n8610), .A1(n8637), .S(n3477), .Z(N2778) );
  CMX2X1 U18050 ( .A0(mem_data1[717]), .A1(mem_data1[718]), .S(n3867), .Z(
        n8617) );
  CMXI2X1 U18051 ( .A0(n8617), .A1(n8611), .S(n4029), .Z(n8624) );
  CMX2X1 U18052 ( .A0(n8612), .A1(n8624), .S(n4342), .Z(n8640) );
  CMXI2X1 U18053 ( .A0(n8613), .A1(n8640), .S(n3477), .Z(N2779) );
  CMX2X1 U18054 ( .A0(mem_data1[718]), .A1(mem_data1[719]), .S(n3875), .Z(
        n8620) );
  CMXI2X1 U18055 ( .A0(n8620), .A1(n8614), .S(n4029), .Z(n8627) );
  CMX2X1 U18056 ( .A0(n8615), .A1(n8627), .S(n4342), .Z(n8643) );
  CMXI2X1 U18057 ( .A0(n8616), .A1(n8643), .S(n3477), .Z(N2780) );
  CMX2X1 U18058 ( .A0(mem_data1[719]), .A1(mem_data1[720]), .S(n3876), .Z(
        n8623) );
  CMXI2X1 U18059 ( .A0(n8623), .A1(n8617), .S(n4029), .Z(n8630) );
  CMX2X1 U18060 ( .A0(n8618), .A1(n8630), .S(n4342), .Z(n8646) );
  CMXI2X1 U18061 ( .A0(n8619), .A1(n8646), .S(n3477), .Z(N2781) );
  CMX2X1 U18062 ( .A0(mem_data1[720]), .A1(mem_data1[721]), .S(n3877), .Z(
        n8626) );
  CMXI2X1 U18063 ( .A0(n8626), .A1(n8620), .S(n4029), .Z(n8636) );
  CMX2X1 U18064 ( .A0(n8621), .A1(n8636), .S(n4342), .Z(n8649) );
  CMXI2X1 U18065 ( .A0(n8622), .A1(n8649), .S(n3477), .Z(N2782) );
  CMX2X1 U18066 ( .A0(mem_data1[721]), .A1(mem_data1[722]), .S(n3878), .Z(
        n8629) );
  CMXI2X1 U18067 ( .A0(n8629), .A1(n8623), .S(n4029), .Z(n8639) );
  CMX2X1 U18068 ( .A0(n8624), .A1(n8639), .S(n4342), .Z(n8652) );
  CMXI2X1 U18069 ( .A0(n8625), .A1(n8652), .S(n3476), .Z(N2783) );
  CMX2X1 U18070 ( .A0(mem_data1[722]), .A1(mem_data1[723]), .S(n3879), .Z(
        n8635) );
  CMXI2X1 U18071 ( .A0(n8635), .A1(n8626), .S(n4029), .Z(n8642) );
  CMX2X1 U18072 ( .A0(n8627), .A1(n8642), .S(n4323), .Z(n8655) );
  CMXI2X1 U18073 ( .A0(n8628), .A1(n8655), .S(n3476), .Z(N2784) );
  CMX2X1 U18074 ( .A0(mem_data1[723]), .A1(mem_data1[724]), .S(n3862), .Z(
        n8638) );
  CMXI2X1 U18075 ( .A0(n8638), .A1(n8629), .S(n4029), .Z(n8645) );
  CMX2X1 U18076 ( .A0(n8630), .A1(n8645), .S(n4369), .Z(n8658) );
  CMXI2X1 U18077 ( .A0(n8631), .A1(n8658), .S(n3476), .Z(N2785) );
  CMX2X1 U18078 ( .A0(mem_data1[84]), .A1(mem_data1[85]), .S(n3863), .Z(n8698)
         );
  CMXI2X1 U18079 ( .A0(n8698), .A1(n8632), .S(n4028), .Z(n8765) );
  CMX2X1 U18080 ( .A0(n8633), .A1(n8765), .S(n4328), .Z(n8898) );
  CMXI2X1 U18081 ( .A0(n8634), .A1(n8898), .S(n3476), .Z(N2146) );
  CMX2X1 U18082 ( .A0(mem_data1[724]), .A1(mem_data1[725]), .S(n3880), .Z(
        n8641) );
  CMXI2X1 U18083 ( .A0(n8641), .A1(n8635), .S(n4028), .Z(n8648) );
  CMX2X1 U18084 ( .A0(n8636), .A1(n8648), .S(n4374), .Z(n8661) );
  CMXI2X1 U18085 ( .A0(n8637), .A1(n8661), .S(n3476), .Z(N2786) );
  CMX2X1 U18086 ( .A0(mem_data1[725]), .A1(mem_data1[726]), .S(n3881), .Z(
        n8644) );
  CMXI2X1 U18087 ( .A0(n8644), .A1(n8638), .S(n4028), .Z(n8651) );
  CMX2X1 U18088 ( .A0(n8639), .A1(n8651), .S(n4373), .Z(n8664) );
  CMXI2X1 U18089 ( .A0(n8640), .A1(n8664), .S(n3476), .Z(N2787) );
  CMX2X1 U18090 ( .A0(mem_data1[726]), .A1(mem_data1[727]), .S(n3868), .Z(
        n8647) );
  CMXI2X1 U18091 ( .A0(n8647), .A1(n8641), .S(n4028), .Z(n8654) );
  CMX2X1 U18092 ( .A0(n8642), .A1(n8654), .S(n4334), .Z(n8670) );
  CMXI2X1 U18093 ( .A0(n8643), .A1(n8670), .S(n3476), .Z(N2788) );
  CMX2X1 U18094 ( .A0(mem_data1[727]), .A1(mem_data1[728]), .S(n3869), .Z(
        n8650) );
  CMXI2X1 U18095 ( .A0(n8650), .A1(n8644), .S(n4028), .Z(n8657) );
  CMX2X1 U18096 ( .A0(n8645), .A1(n8657), .S(n4335), .Z(n8673) );
  CMXI2X1 U18097 ( .A0(n8646), .A1(n8673), .S(n3476), .Z(N2789) );
  CMX2X1 U18098 ( .A0(mem_data1[728]), .A1(mem_data1[729]), .S(n3870), .Z(
        n8653) );
  CMXI2X1 U18099 ( .A0(n8653), .A1(n8647), .S(n4028), .Z(n8660) );
  CMX2X1 U18100 ( .A0(n8648), .A1(n8660), .S(n4324), .Z(n8676) );
  CMXI2X1 U18101 ( .A0(n8649), .A1(n8676), .S(n3476), .Z(N2790) );
  CMX2X1 U18102 ( .A0(mem_data1[729]), .A1(mem_data1[730]), .S(n3871), .Z(
        n8656) );
  CMXI2X1 U18103 ( .A0(n8656), .A1(n8650), .S(n4028), .Z(n8663) );
  CMX2X1 U18104 ( .A0(n8651), .A1(n8663), .S(n4325), .Z(n8679) );
  CMXI2X1 U18105 ( .A0(n8652), .A1(n8679), .S(n3479), .Z(N2791) );
  CMX2X1 U18106 ( .A0(mem_data1[730]), .A1(mem_data1[731]), .S(n3868), .Z(
        n8659) );
  CMXI2X1 U18107 ( .A0(n8659), .A1(n8653), .S(n4028), .Z(n8669) );
  CMX2X1 U18108 ( .A0(n8654), .A1(n8669), .S(n4326), .Z(n8682) );
  CMXI2X1 U18109 ( .A0(n8655), .A1(n8682), .S(n3479), .Z(N2792) );
  CMX2X1 U18110 ( .A0(mem_data1[731]), .A1(mem_data1[732]), .S(n3869), .Z(
        n8662) );
  CMXI2X1 U18111 ( .A0(n8662), .A1(n8656), .S(n4028), .Z(n8672) );
  CMX2X1 U18112 ( .A0(n8657), .A1(n8672), .S(n4327), .Z(n8685) );
  CMXI2X1 U18113 ( .A0(n8658), .A1(n8685), .S(n3479), .Z(N2793) );
  CMX2X1 U18114 ( .A0(mem_data1[732]), .A1(mem_data1[733]), .S(n3870), .Z(
        n8668) );
  CMXI2X1 U18115 ( .A0(n8668), .A1(n8659), .S(n4028), .Z(n8675) );
  CMX2X1 U18116 ( .A0(n8660), .A1(n8675), .S(n4341), .Z(n8688) );
  CMXI2X1 U18117 ( .A0(n8661), .A1(n8688), .S(n3479), .Z(N2794) );
  CMX2X1 U18118 ( .A0(mem_data1[733]), .A1(mem_data1[734]), .S(n3871), .Z(
        n8671) );
  CMXI2X1 U18119 ( .A0(n8671), .A1(n8662), .S(n4028), .Z(n8678) );
  CMX2X1 U18120 ( .A0(n8663), .A1(n8678), .S(n4341), .Z(n8691) );
  CMXI2X1 U18121 ( .A0(n8664), .A1(n8691), .S(n3479), .Z(N2795) );
  CMX2X1 U18122 ( .A0(mem_data1[85]), .A1(mem_data1[86]), .S(n3873), .Z(n8731)
         );
  CMXI2X1 U18123 ( .A0(n8731), .A1(n8665), .S(n4028), .Z(n8798) );
  CMX2X1 U18124 ( .A0(n8666), .A1(n8798), .S(n4341), .Z(n8931) );
  CMXI2X1 U18125 ( .A0(n8667), .A1(n8931), .S(n3478), .Z(N2147) );
  CMX2X1 U18126 ( .A0(mem_data1[734]), .A1(mem_data1[735]), .S(n3862), .Z(
        n8674) );
  CMXI2X1 U18127 ( .A0(n8674), .A1(n8668), .S(n4028), .Z(n8681) );
  CMX2X1 U18128 ( .A0(n8669), .A1(n8681), .S(n4341), .Z(n8694) );
  CMXI2X1 U18129 ( .A0(n8670), .A1(n8694), .S(n3478), .Z(N2796) );
  CMX2X1 U18130 ( .A0(mem_data1[735]), .A1(mem_data1[736]), .S(n3863), .Z(
        n8677) );
  CMXI2X1 U18131 ( .A0(n8677), .A1(n8671), .S(n4028), .Z(n8684) );
  CMX2X1 U18132 ( .A0(n8672), .A1(n8684), .S(n4341), .Z(n8697) );
  CMXI2X1 U18133 ( .A0(n8673), .A1(n8697), .S(n3478), .Z(N2797) );
  CMX2X1 U18134 ( .A0(mem_data1[736]), .A1(mem_data1[737]), .S(n3864), .Z(
        n8680) );
  CMXI2X1 U18135 ( .A0(n8680), .A1(n8674), .S(n4028), .Z(n8687) );
  CMX2X1 U18136 ( .A0(n8675), .A1(n8687), .S(n4341), .Z(n8703) );
  CMXI2X1 U18137 ( .A0(n8676), .A1(n8703), .S(n3478), .Z(N2798) );
  CMX2X1 U18138 ( .A0(mem_data1[737]), .A1(mem_data1[738]), .S(n3865), .Z(
        n8683) );
  CMXI2X1 U18139 ( .A0(n8683), .A1(n8677), .S(n4028), .Z(n8690) );
  CMX2X1 U18140 ( .A0(n8678), .A1(n8690), .S(n4341), .Z(n8706) );
  CMXI2X1 U18141 ( .A0(n8679), .A1(n8706), .S(n3478), .Z(N2799) );
  CMX2X1 U18142 ( .A0(mem_data1[738]), .A1(mem_data1[739]), .S(n3866), .Z(
        n8686) );
  CMXI2X1 U18143 ( .A0(n8686), .A1(n8680), .S(n4027), .Z(n8693) );
  CMX2X1 U18144 ( .A0(n8681), .A1(n8693), .S(n4341), .Z(n8709) );
  CMXI2X1 U18145 ( .A0(n8682), .A1(n8709), .S(n3478), .Z(N2800) );
  CMX2X1 U18146 ( .A0(mem_data1[739]), .A1(mem_data1[740]), .S(n3867), .Z(
        n8689) );
  CMXI2X1 U18147 ( .A0(n8689), .A1(n8683), .S(n4027), .Z(n8696) );
  CMX2X1 U18148 ( .A0(n8684), .A1(n8696), .S(n4341), .Z(n8712) );
  CMXI2X1 U18149 ( .A0(n8685), .A1(n8712), .S(n3478), .Z(N2801) );
  CMX2X1 U18150 ( .A0(mem_data1[740]), .A1(mem_data1[741]), .S(n3872), .Z(
        n8692) );
  CMXI2X1 U18151 ( .A0(n8692), .A1(n8686), .S(n4027), .Z(n8702) );
  CMX2X1 U18152 ( .A0(n8687), .A1(n8702), .S(n4341), .Z(n8715) );
  CMXI2X1 U18153 ( .A0(n8688), .A1(n8715), .S(n3478), .Z(N2802) );
  CMX2X1 U18154 ( .A0(mem_data1[741]), .A1(mem_data1[742]), .S(n3873), .Z(
        n8695) );
  CMXI2X1 U18155 ( .A0(n8695), .A1(n8689), .S(n4027), .Z(n8705) );
  CMX2X1 U18156 ( .A0(n8690), .A1(n8705), .S(n4341), .Z(n8718) );
  CMXI2X1 U18157 ( .A0(n8691), .A1(n8718), .S(n3478), .Z(N2803) );
  CMX2X1 U18158 ( .A0(mem_data1[742]), .A1(mem_data1[743]), .S(n3874), .Z(
        n8701) );
  CMXI2X1 U18159 ( .A0(n8701), .A1(n8692), .S(n4027), .Z(n8708) );
  CMX2X1 U18160 ( .A0(n8693), .A1(n8708), .S(n4340), .Z(n8721) );
  CMXI2X1 U18161 ( .A0(n8694), .A1(n8721), .S(n3478), .Z(N2804) );
  CMX2X1 U18162 ( .A0(mem_data1[743]), .A1(mem_data1[744]), .S(n3875), .Z(
        n8704) );
  CMXI2X1 U18163 ( .A0(n8704), .A1(n8695), .S(n4027), .Z(n8711) );
  CMX2X1 U18164 ( .A0(n8696), .A1(n8711), .S(n4340), .Z(n8724) );
  CMXI2X1 U18165 ( .A0(n8697), .A1(n8724), .S(n3478), .Z(N2805) );
  CMX2X1 U18166 ( .A0(mem_data1[86]), .A1(mem_data1[87]), .S(n3865), .Z(n8764)
         );
  CMXI2X1 U18167 ( .A0(n8764), .A1(n8698), .S(n4027), .Z(n8831) );
  CMX2X1 U18168 ( .A0(n8699), .A1(n8831), .S(n4340), .Z(n8968) );
  CMXI2X1 U18169 ( .A0(n8700), .A1(n8968), .S(n3477), .Z(N2148) );
  CMX2X1 U18170 ( .A0(mem_data1[744]), .A1(mem_data1[745]), .S(n3866), .Z(
        n8707) );
  CMXI2X1 U18171 ( .A0(n8707), .A1(n8701), .S(n4027), .Z(n8714) );
  CMX2X1 U18172 ( .A0(n8702), .A1(n8714), .S(n4340), .Z(n8727) );
  CMXI2X1 U18173 ( .A0(n8703), .A1(n8727), .S(n3477), .Z(N2806) );
  CMX2X1 U18174 ( .A0(mem_data1[745]), .A1(mem_data1[746]), .S(n3867), .Z(
        n8710) );
  CMXI2X1 U18175 ( .A0(n8710), .A1(n8704), .S(n4027), .Z(n8717) );
  CMX2X1 U18176 ( .A0(n8705), .A1(n8717), .S(n4340), .Z(n8730) );
  CMXI2X1 U18177 ( .A0(n8706), .A1(n8730), .S(n3481), .Z(N2807) );
  CMX2X1 U18178 ( .A0(mem_data1[746]), .A1(mem_data1[747]), .S(n3868), .Z(
        n8713) );
  CMXI2X1 U18179 ( .A0(n8713), .A1(n8707), .S(n4027), .Z(n8720) );
  CMX2X1 U18180 ( .A0(n8708), .A1(n8720), .S(n4340), .Z(n8736) );
  CMXI2X1 U18181 ( .A0(n8709), .A1(n8736), .S(n3480), .Z(N2808) );
  CMX2X1 U18182 ( .A0(mem_data1[747]), .A1(mem_data1[748]), .S(n3864), .Z(
        n8716) );
  CMXI2X1 U18183 ( .A0(n8716), .A1(n8710), .S(n4027), .Z(n8723) );
  CMX2X1 U18184 ( .A0(n8711), .A1(n8723), .S(n4340), .Z(n8739) );
  CMXI2X1 U18185 ( .A0(n8712), .A1(n8739), .S(n3480), .Z(N2809) );
  CMX2X1 U18186 ( .A0(mem_data1[748]), .A1(mem_data1[749]), .S(n3868), .Z(
        n8719) );
  CMXI2X1 U18187 ( .A0(n8719), .A1(n8713), .S(n4027), .Z(n8726) );
  CMX2X1 U18188 ( .A0(n8714), .A1(n8726), .S(n4340), .Z(n8742) );
  CMXI2X1 U18189 ( .A0(n8715), .A1(n8742), .S(n3480), .Z(N2810) );
  CMX2X1 U18190 ( .A0(mem_data1[749]), .A1(mem_data1[750]), .S(n3869), .Z(
        n8722) );
  CMXI2X1 U18191 ( .A0(n8722), .A1(n8716), .S(n4027), .Z(n8729) );
  CMX2X1 U18192 ( .A0(n8717), .A1(n8729), .S(n4340), .Z(n8745) );
  CMXI2X1 U18193 ( .A0(n8718), .A1(n8745), .S(n3480), .Z(N2811) );
  CMX2X1 U18194 ( .A0(mem_data1[750]), .A1(mem_data1[751]), .S(n3870), .Z(
        n8725) );
  CMXI2X1 U18195 ( .A0(n8725), .A1(n8719), .S(n4027), .Z(n8735) );
  CMX2X1 U18196 ( .A0(n8720), .A1(n8735), .S(n4340), .Z(n8748) );
  CMXI2X1 U18197 ( .A0(n8721), .A1(n8748), .S(n3480), .Z(N2812) );
  CMX2X1 U18198 ( .A0(mem_data1[751]), .A1(mem_data1[752]), .S(n3871), .Z(
        n8728) );
  CMXI2X1 U18199 ( .A0(n8728), .A1(n8722), .S(n4027), .Z(n8738) );
  CMX2X1 U18200 ( .A0(n8723), .A1(n8738), .S(n4340), .Z(n8751) );
  CMXI2X1 U18201 ( .A0(n8724), .A1(n8751), .S(n3480), .Z(N2813) );
  CMX2X1 U18202 ( .A0(mem_data1[752]), .A1(mem_data1[753]), .S(n3872), .Z(
        n8734) );
  CMXI2X1 U18203 ( .A0(n8734), .A1(n8725), .S(n4027), .Z(n8741) );
  CMX2X1 U18204 ( .A0(n8726), .A1(n8741), .S(n4340), .Z(n8754) );
  CMXI2X1 U18205 ( .A0(n8727), .A1(n8754), .S(n3480), .Z(N2814) );
  CMX2X1 U18206 ( .A0(mem_data1[753]), .A1(mem_data1[754]), .S(n3873), .Z(
        n8737) );
  CMXI2X1 U18207 ( .A0(n8737), .A1(n8728), .S(n4026), .Z(n8744) );
  CMX2X1 U18208 ( .A0(n8729), .A1(n8744), .S(n4338), .Z(n8757) );
  CMXI2X1 U18209 ( .A0(n8730), .A1(n8757), .S(n3480), .Z(N2815) );
  CMX2X1 U18210 ( .A0(mem_data1[87]), .A1(mem_data1[88]), .S(n3874), .Z(n8797)
         );
  CMXI2X1 U18211 ( .A0(n8797), .A1(n8731), .S(n4026), .Z(n8864) );
  CMX2X1 U18212 ( .A0(n8732), .A1(n8864), .S(n4365), .Z(n9001) );
  CMXI2X1 U18213 ( .A0(n8733), .A1(n9001), .S(n3480), .Z(N2149) );
  CMX2X1 U18214 ( .A0(mem_data1[754]), .A1(mem_data1[755]), .S(n3868), .Z(
        n8740) );
  CMXI2X1 U18215 ( .A0(n8740), .A1(n8734), .S(n4026), .Z(n8747) );
  CMX2X1 U18216 ( .A0(n8735), .A1(n8747), .S(n4329), .Z(n8760) );
  CMXI2X1 U18217 ( .A0(n8736), .A1(n8760), .S(n3480), .Z(N2816) );
  CMX2X1 U18218 ( .A0(mem_data1[755]), .A1(mem_data1[756]), .S(n3869), .Z(
        n8743) );
  CMXI2X1 U18219 ( .A0(n8743), .A1(n8737), .S(n4026), .Z(n8750) );
  CMX2X1 U18220 ( .A0(n8738), .A1(n8750), .S(n4330), .Z(n8763) );
  CMXI2X1 U18221 ( .A0(n8739), .A1(n8763), .S(n3480), .Z(N2817) );
  CMX2X1 U18222 ( .A0(mem_data1[756]), .A1(mem_data1[757]), .S(n3875), .Z(
        n8746) );
  CMXI2X1 U18223 ( .A0(n8746), .A1(n8740), .S(n4026), .Z(n8753) );
  CMX2X1 U18224 ( .A0(n8741), .A1(n8753), .S(n4323), .Z(n8769) );
  CMXI2X1 U18225 ( .A0(n8742), .A1(n8769), .S(n3479), .Z(N2818) );
  CMX2X1 U18226 ( .A0(mem_data1[757]), .A1(mem_data1[758]), .S(n3875), .Z(
        n8749) );
  CMXI2X1 U18227 ( .A0(n8749), .A1(n8743), .S(n4026), .Z(n8756) );
  CMX2X1 U18228 ( .A0(n8744), .A1(n8756), .S(n4325), .Z(n8772) );
  CMXI2X1 U18229 ( .A0(n8745), .A1(n8772), .S(n3479), .Z(N2819) );
  CMX2X1 U18230 ( .A0(mem_data1[758]), .A1(mem_data1[759]), .S(n3869), .Z(
        n8752) );
  CMXI2X1 U18231 ( .A0(n8752), .A1(n8746), .S(n4026), .Z(n8759) );
  CMX2X1 U18232 ( .A0(n8747), .A1(n8759), .S(n4328), .Z(n8775) );
  CMXI2X1 U18233 ( .A0(n8748), .A1(n8775), .S(n3479), .Z(N2820) );
  CMX2X1 U18234 ( .A0(mem_data1[759]), .A1(mem_data1[760]), .S(n4278), .Z(
        n8755) );
  CMXI2X1 U18235 ( .A0(n8755), .A1(n8749), .S(n4026), .Z(n8762) );
  CMX2X1 U18236 ( .A0(n8750), .A1(n8762), .S(n4372), .Z(n8778) );
  CMXI2X1 U18237 ( .A0(n8751), .A1(n8778), .S(n3479), .Z(N2821) );
  CMX2X1 U18238 ( .A0(mem_data1[760]), .A1(mem_data1[761]), .S(n4278), .Z(
        n8758) );
  CMXI2X1 U18239 ( .A0(n8758), .A1(n8752), .S(n4026), .Z(n8768) );
  CMX2X1 U18240 ( .A0(n8753), .A1(n8768), .S(n4368), .Z(n8781) );
  CMXI2X1 U18241 ( .A0(n8754), .A1(n8781), .S(n3479), .Z(N2822) );
  CMX2X1 U18242 ( .A0(mem_data1[761]), .A1(mem_data1[762]), .S(n4278), .Z(
        n8761) );
  CMXI2X1 U18243 ( .A0(n8761), .A1(n8755), .S(n4026), .Z(n8771) );
  CMX2X1 U18244 ( .A0(n8756), .A1(n8771), .S(n4375), .Z(n8784) );
  CMXI2X1 U18245 ( .A0(n8757), .A1(n8784), .S(n3479), .Z(N2823) );
  CMX2X1 U18246 ( .A0(mem_data1[762]), .A1(mem_data1[763]), .S(n4278), .Z(
        n8767) );
  CMXI2X1 U18247 ( .A0(n8767), .A1(n8758), .S(n4026), .Z(n8774) );
  CMX2X1 U18248 ( .A0(n8759), .A1(n8774), .S(n4339), .Z(n8787) );
  CMXI2X1 U18249 ( .A0(n8760), .A1(n8787), .S(n3517), .Z(N2824) );
  CMX2X1 U18250 ( .A0(mem_data1[763]), .A1(mem_data1[764]), .S(n4278), .Z(
        n8770) );
  CMXI2X1 U18251 ( .A0(n8770), .A1(n8761), .S(n4026), .Z(n8777) );
  CMX2X1 U18252 ( .A0(n8762), .A1(n8777), .S(n4339), .Z(n8790) );
  CMXI2X1 U18253 ( .A0(n8763), .A1(n8790), .S(n3517), .Z(N2825) );
  CMX2X1 U18254 ( .A0(mem_data1[88]), .A1(mem_data1[89]), .S(n4278), .Z(n8830)
         );
  CMXI2X1 U18255 ( .A0(n8830), .A1(n8764), .S(n4026), .Z(n8897) );
  CMX2X1 U18256 ( .A0(n8765), .A1(n8897), .S(n4339), .Z(n9034) );
  CMXI2X1 U18257 ( .A0(n8766), .A1(n9034), .S(n3517), .Z(N2150) );
  CMX2X1 U18258 ( .A0(mem_data1[764]), .A1(mem_data1[765]), .S(n4278), .Z(
        n8773) );
  CMXI2X1 U18259 ( .A0(n8773), .A1(n8767), .S(n4026), .Z(n8780) );
  CMX2X1 U18260 ( .A0(n8768), .A1(n8780), .S(n4339), .Z(n8793) );
  CMXI2X1 U18261 ( .A0(n8769), .A1(n8793), .S(n3517), .Z(N2826) );
  CMX2X1 U18262 ( .A0(mem_data1[765]), .A1(mem_data1[766]), .S(n4277), .Z(
        n8776) );
  CMXI2X1 U18263 ( .A0(n8776), .A1(n8770), .S(n4026), .Z(n8783) );
  CMX2X1 U18264 ( .A0(n8771), .A1(n8783), .S(n4339), .Z(n8796) );
  CMXI2X1 U18265 ( .A0(n8772), .A1(n8796), .S(n3516), .Z(N2827) );
  CMX2X1 U18266 ( .A0(mem_data1[766]), .A1(mem_data1[767]), .S(n4277), .Z(
        n8779) );
  CMXI2X1 U18267 ( .A0(n8779), .A1(n8773), .S(n4026), .Z(n8786) );
  CMX2X1 U18268 ( .A0(n8774), .A1(n8786), .S(n4339), .Z(n8802) );
  CMXI2X1 U18269 ( .A0(n8775), .A1(n8802), .S(n3516), .Z(N2828) );
  CMX2X1 U18270 ( .A0(mem_data1[767]), .A1(mem_data1[768]), .S(n4277), .Z(
        n8782) );
  CMXI2X1 U18271 ( .A0(n8782), .A1(n8776), .S(n4025), .Z(n8789) );
  CMX2X1 U18272 ( .A0(n8777), .A1(n8789), .S(n4339), .Z(n8805) );
  CMXI2X1 U18273 ( .A0(n8778), .A1(n8805), .S(n3516), .Z(N2829) );
  CMX2X1 U18274 ( .A0(mem_data1[768]), .A1(mem_data1[769]), .S(n4277), .Z(
        n8785) );
  CMXI2X1 U18275 ( .A0(n8785), .A1(n8779), .S(n4025), .Z(n8792) );
  CMX2X1 U18276 ( .A0(n8780), .A1(n8792), .S(n4342), .Z(n8808) );
  CMXI2X1 U18277 ( .A0(n8781), .A1(n8808), .S(n3349), .Z(N2830) );
  CMX2X1 U18278 ( .A0(mem_data1[769]), .A1(mem_data1[770]), .S(n4277), .Z(
        n8788) );
  CMXI2X1 U18279 ( .A0(n8788), .A1(n8782), .S(n4025), .Z(n8795) );
  CMX2X1 U18280 ( .A0(n8783), .A1(n8795), .S(n4353), .Z(n8811) );
  CMXI2X1 U18281 ( .A0(n8784), .A1(n8811), .S(n3516), .Z(N2831) );
  CMX2X1 U18282 ( .A0(mem_data1[770]), .A1(mem_data1[771]), .S(n4277), .Z(
        n8791) );
  CMXI2X1 U18283 ( .A0(n8791), .A1(n8785), .S(n4025), .Z(n8801) );
  CMX2X1 U18284 ( .A0(n8786), .A1(n8801), .S(n3808), .Z(n8814) );
  CMXI2X1 U18285 ( .A0(n8787), .A1(n8814), .S(n3516), .Z(N2832) );
  CMX2X1 U18286 ( .A0(mem_data1[771]), .A1(mem_data1[772]), .S(n4277), .Z(
        n8794) );
  CMXI2X1 U18287 ( .A0(n8794), .A1(n8788), .S(n4025), .Z(n8804) );
  CMX2X1 U18288 ( .A0(n8789), .A1(n8804), .S(n3809), .Z(n8817) );
  CMXI2X1 U18289 ( .A0(n8790), .A1(n8817), .S(n3516), .Z(N2833) );
  CMX2X1 U18290 ( .A0(mem_data1[772]), .A1(mem_data1[773]), .S(n4277), .Z(
        n8800) );
  CMXI2X1 U18291 ( .A0(n8800), .A1(n8791), .S(n4025), .Z(n8807) );
  CMX2X1 U18292 ( .A0(n8792), .A1(n8807), .S(n3810), .Z(n8820) );
  CMXI2X1 U18293 ( .A0(n8793), .A1(n8820), .S(n3516), .Z(N2834) );
  CMX2X1 U18294 ( .A0(mem_data1[773]), .A1(mem_data1[774]), .S(n4277), .Z(
        n8803) );
  CMXI2X1 U18295 ( .A0(n8803), .A1(n8794), .S(n4025), .Z(n8810) );
  CMX2X1 U18296 ( .A0(n8795), .A1(n8810), .S(n3811), .Z(n8823) );
  CMXI2X1 U18297 ( .A0(n8796), .A1(n8823), .S(n3516), .Z(N2835) );
  CMX2X1 U18298 ( .A0(mem_data1[89]), .A1(mem_data1[90]), .S(n4277), .Z(n8863)
         );
  CMXI2X1 U18299 ( .A0(n8863), .A1(n8797), .S(n4025), .Z(n8930) );
  CMX2X1 U18300 ( .A0(n8798), .A1(n8930), .S(n3794), .Z(n9067) );
  CMXI2X1 U18301 ( .A0(n8799), .A1(n9067), .S(n3516), .Z(N2151) );
  CMX2X1 U18302 ( .A0(mem_data1[774]), .A1(mem_data1[775]), .S(n4277), .Z(
        n8806) );
  CMXI2X1 U18303 ( .A0(n8806), .A1(n8800), .S(n4025), .Z(n8813) );
  CMX2X1 U18304 ( .A0(n8801), .A1(n8813), .S(n3807), .Z(n8826) );
  CMXI2X1 U18305 ( .A0(n8802), .A1(n8826), .S(n3516), .Z(N2836) );
  CMX2X1 U18306 ( .A0(mem_data1[775]), .A1(mem_data1[776]), .S(n4276), .Z(
        n8809) );
  CMXI2X1 U18307 ( .A0(n8809), .A1(n8803), .S(n4025), .Z(n8816) );
  CMX2X1 U18308 ( .A0(n8804), .A1(n8816), .S(n3808), .Z(n8829) );
  CMXI2X1 U18309 ( .A0(n8805), .A1(n8829), .S(n3516), .Z(N2837) );
  CMX2X1 U18310 ( .A0(mem_data1[776]), .A1(mem_data1[777]), .S(n4276), .Z(
        n8812) );
  CMXI2X1 U18311 ( .A0(n8812), .A1(n8806), .S(n4025), .Z(n8819) );
  CMX2X1 U18312 ( .A0(n8807), .A1(n8819), .S(n3809), .Z(n8835) );
  CMXI2X1 U18313 ( .A0(n8808), .A1(n8835), .S(n3515), .Z(N2838) );
  CMX2X1 U18314 ( .A0(mem_data1[777]), .A1(mem_data1[778]), .S(n4276), .Z(
        n8815) );
  CMXI2X1 U18315 ( .A0(n8815), .A1(n8809), .S(n4025), .Z(n8822) );
  CMX2X1 U18316 ( .A0(n8810), .A1(n8822), .S(n3810), .Z(n8838) );
  CMXI2X1 U18317 ( .A0(n8811), .A1(n8838), .S(n3515), .Z(N2839) );
  CMX2X1 U18318 ( .A0(mem_data1[778]), .A1(mem_data1[779]), .S(n4276), .Z(
        n8818) );
  CMXI2X1 U18319 ( .A0(n8818), .A1(n8812), .S(n4025), .Z(n8825) );
  CMX2X1 U18320 ( .A0(n8813), .A1(n8825), .S(n3811), .Z(n8841) );
  CMXI2X1 U18321 ( .A0(n8814), .A1(n8841), .S(n3517), .Z(N2840) );
  CMX2X1 U18322 ( .A0(mem_data1[779]), .A1(mem_data1[780]), .S(n4276), .Z(
        n8821) );
  CMXI2X1 U18323 ( .A0(n8821), .A1(n8815), .S(n4025), .Z(n8828) );
  CMX2X1 U18324 ( .A0(n8816), .A1(n8828), .S(n3812), .Z(n8844) );
  CMXI2X1 U18325 ( .A0(n8817), .A1(n8844), .S(n3518), .Z(N2841) );
  CMX2X1 U18326 ( .A0(mem_data1[780]), .A1(mem_data1[781]), .S(n4276), .Z(
        n8824) );
  CMXI2X1 U18327 ( .A0(n8824), .A1(n8818), .S(n4025), .Z(n8834) );
  CMX2X1 U18328 ( .A0(n8819), .A1(n8834), .S(n4356), .Z(n8847) );
  CMXI2X1 U18329 ( .A0(n8820), .A1(n8847), .S(n3518), .Z(N2842) );
  CMX2X1 U18330 ( .A0(mem_data1[781]), .A1(mem_data1[782]), .S(n4276), .Z(
        n8827) );
  CMXI2X1 U18331 ( .A0(n8827), .A1(n8821), .S(n4025), .Z(n8837) );
  CMX2X1 U18332 ( .A0(n8822), .A1(n8837), .S(n3771), .Z(n8850) );
  CMXI2X1 U18333 ( .A0(n8823), .A1(n8850), .S(n3518), .Z(N2843) );
  CMX2X1 U18334 ( .A0(mem_data1[782]), .A1(mem_data1[783]), .S(n4276), .Z(
        n8833) );
  CMXI2X1 U18335 ( .A0(n8833), .A1(n8824), .S(n4024), .Z(n8840) );
  CMX2X1 U18336 ( .A0(n8825), .A1(n8840), .S(n3772), .Z(n8853) );
  CMXI2X1 U18337 ( .A0(n8826), .A1(n8853), .S(n3471), .Z(N2844) );
  CMX2X1 U18338 ( .A0(mem_data1[783]), .A1(mem_data1[784]), .S(n4276), .Z(
        n8836) );
  CMXI2X1 U18339 ( .A0(n8836), .A1(n8827), .S(n4024), .Z(n8843) );
  CMX2X1 U18340 ( .A0(n8828), .A1(n8843), .S(n3773), .Z(n8856) );
  CMXI2X1 U18341 ( .A0(n8829), .A1(n8856), .S(n3325), .Z(N2845) );
  CMX2X1 U18342 ( .A0(mem_data1[90]), .A1(mem_data1[91]), .S(n4276), .Z(n8896)
         );
  CMXI2X1 U18343 ( .A0(n8896), .A1(n8830), .S(n4024), .Z(n8967) );
  CMX2X1 U18344 ( .A0(n8831), .A1(n8967), .S(n3774), .Z(n9100) );
  CMXI2X1 U18345 ( .A0(n8832), .A1(n9100), .S(n3317), .Z(N2152) );
  CMX2X1 U18346 ( .A0(mem_data1[784]), .A1(mem_data1[785]), .S(n4276), .Z(
        n8839) );
  CMXI2X1 U18347 ( .A0(n8839), .A1(n8833), .S(n4024), .Z(n8846) );
  CMX2X1 U18348 ( .A0(n8834), .A1(n8846), .S(n3775), .Z(n8859) );
  CMXI2X1 U18349 ( .A0(n8835), .A1(n8859), .S(n3317), .Z(N2846) );
  CMX2X1 U18350 ( .A0(mem_data1[785]), .A1(mem_data1[786]), .S(n4275), .Z(
        n8842) );
  CMXI2X1 U18351 ( .A0(n8842), .A1(n8836), .S(n4024), .Z(n8849) );
  CMX2X1 U18352 ( .A0(n8837), .A1(n8849), .S(n3776), .Z(n8862) );
  CMXI2X1 U18353 ( .A0(n8838), .A1(n8862), .S(n3316), .Z(N2847) );
  CMX2X1 U18354 ( .A0(mem_data1[786]), .A1(mem_data1[787]), .S(n4275), .Z(
        n8845) );
  CMXI2X1 U18355 ( .A0(n8845), .A1(n8839), .S(n4024), .Z(n8852) );
  CMX2X1 U18356 ( .A0(n8840), .A1(n8852), .S(n3777), .Z(n8868) );
  CMXI2X1 U18357 ( .A0(n8841), .A1(n8868), .S(n3316), .Z(N2848) );
  CMX2X1 U18358 ( .A0(mem_data1[787]), .A1(mem_data1[788]), .S(n4275), .Z(
        n8848) );
  CMXI2X1 U18359 ( .A0(n8848), .A1(n8842), .S(n4024), .Z(n8855) );
  CMX2X1 U18360 ( .A0(n8843), .A1(n8855), .S(n3790), .Z(n8871) );
  CMXI2X1 U18361 ( .A0(n8844), .A1(n8871), .S(n3316), .Z(N2849) );
  CMX2X1 U18362 ( .A0(mem_data1[788]), .A1(mem_data1[789]), .S(n4275), .Z(
        n8851) );
  CMXI2X1 U18363 ( .A0(n8851), .A1(n8845), .S(n4024), .Z(n8858) );
  CMX2X1 U18364 ( .A0(n8846), .A1(n8858), .S(n3791), .Z(n8874) );
  CMXI2X1 U18365 ( .A0(n8847), .A1(n8874), .S(n3316), .Z(N2850) );
  CMX2X1 U18366 ( .A0(mem_data1[789]), .A1(mem_data1[790]), .S(n4275), .Z(
        n8854) );
  CMXI2X1 U18367 ( .A0(n8854), .A1(n8848), .S(n4024), .Z(n8861) );
  CMX2X1 U18368 ( .A0(n8849), .A1(n8861), .S(n3772), .Z(n8877) );
  CMXI2X1 U18369 ( .A0(n8850), .A1(n8877), .S(n3316), .Z(N2851) );
  CMX2X1 U18370 ( .A0(mem_data1[790]), .A1(mem_data1[791]), .S(n4275), .Z(
        n8857) );
  CMXI2X1 U18371 ( .A0(n8857), .A1(n8851), .S(n4024), .Z(n8867) );
  CMX2X1 U18372 ( .A0(n8852), .A1(n8867), .S(n3771), .Z(n8880) );
  CMXI2X1 U18373 ( .A0(n8853), .A1(n8880), .S(n3316), .Z(N2852) );
  CMX2X1 U18374 ( .A0(mem_data1[791]), .A1(mem_data1[792]), .S(n4275), .Z(
        n8860) );
  CMXI2X1 U18375 ( .A0(n8860), .A1(n8854), .S(n4024), .Z(n8870) );
  CMX2X1 U18376 ( .A0(n8855), .A1(n8870), .S(n3812), .Z(n8883) );
  CMXI2X1 U18377 ( .A0(n8856), .A1(n8883), .S(n3316), .Z(N2853) );
  CMX2X1 U18378 ( .A0(mem_data1[792]), .A1(mem_data1[793]), .S(n4275), .Z(
        n8866) );
  CMXI2X1 U18379 ( .A0(n8866), .A1(n8857), .S(n4024), .Z(n8873) );
  CMX2X1 U18380 ( .A0(n8858), .A1(n8873), .S(n4354), .Z(n8886) );
  CMXI2X1 U18381 ( .A0(n8859), .A1(n8886), .S(n3316), .Z(N2854) );
  CMX2X1 U18382 ( .A0(mem_data1[793]), .A1(mem_data1[794]), .S(n4275), .Z(
        n8869) );
  CMXI2X1 U18383 ( .A0(n8869), .A1(n8860), .S(n4024), .Z(n8876) );
  CMX2X1 U18384 ( .A0(n8861), .A1(n8876), .S(n3771), .Z(n8889) );
  CMXI2X1 U18385 ( .A0(n8862), .A1(n8889), .S(n3316), .Z(N2855) );
  CMX2X1 U18386 ( .A0(mem_data1[91]), .A1(mem_data1[92]), .S(n4275), .Z(n8929)
         );
  CMXI2X1 U18387 ( .A0(n8929), .A1(n8863), .S(n4024), .Z(n9000) );
  CMX2X1 U18388 ( .A0(n8864), .A1(n9000), .S(n3772), .Z(n9133) );
  CMXI2X1 U18389 ( .A0(n8865), .A1(n9133), .S(n3316), .Z(N2153) );
  CMX2X1 U18390 ( .A0(mem_data1[794]), .A1(mem_data1[795]), .S(n4275), .Z(
        n8872) );
  CMXI2X1 U18391 ( .A0(n8872), .A1(n8866), .S(n4024), .Z(n8879) );
  CMX2X1 U18392 ( .A0(n8867), .A1(n8879), .S(n3773), .Z(n8892) );
  CMXI2X1 U18393 ( .A0(n8868), .A1(n8892), .S(n3316), .Z(N2856) );
  CMX2X1 U18394 ( .A0(mem_data1[795]), .A1(mem_data1[796]), .S(n4274), .Z(
        n8875) );
  CMXI2X1 U18395 ( .A0(n8875), .A1(n8869), .S(n4024), .Z(n8882) );
  CMX2X1 U18396 ( .A0(n8870), .A1(n8882), .S(n3795), .Z(n8895) );
  CMXI2X1 U18397 ( .A0(n8871), .A1(n8895), .S(n3315), .Z(N2857) );
  CMX2X1 U18398 ( .A0(mem_data1[796]), .A1(mem_data1[797]), .S(n4274), .Z(
        n8878) );
  CMXI2X1 U18399 ( .A0(n8878), .A1(n8872), .S(n4023), .Z(n8885) );
  CMX2X1 U18400 ( .A0(n8873), .A1(n8885), .S(n3792), .Z(n8901) );
  CMXI2X1 U18401 ( .A0(n8874), .A1(n8901), .S(n3315), .Z(N2858) );
  CMX2X1 U18402 ( .A0(mem_data1[797]), .A1(mem_data1[798]), .S(n4274), .Z(
        n8881) );
  CMXI2X1 U18403 ( .A0(n8881), .A1(n8875), .S(n4023), .Z(n8888) );
  CMX2X1 U18404 ( .A0(n8876), .A1(n8888), .S(n3793), .Z(n8904) );
  CMXI2X1 U18405 ( .A0(n8877), .A1(n8904), .S(n3319), .Z(N2859) );
  CMX2X1 U18406 ( .A0(mem_data1[798]), .A1(mem_data1[799]), .S(n4274), .Z(
        n8884) );
  CMXI2X1 U18407 ( .A0(n8884), .A1(n8878), .S(n4023), .Z(n8891) );
  CMX2X1 U18408 ( .A0(n8879), .A1(n8891), .S(n3794), .Z(n8907) );
  CMXI2X1 U18409 ( .A0(n8880), .A1(n8907), .S(n3318), .Z(N2860) );
  CMX2X1 U18410 ( .A0(mem_data1[799]), .A1(mem_data1[800]), .S(n4274), .Z(
        n8887) );
  CMXI2X1 U18411 ( .A0(n8887), .A1(n8881), .S(n4023), .Z(n8894) );
  CMX2X1 U18412 ( .A0(n8882), .A1(n8894), .S(n3795), .Z(n8910) );
  CMXI2X1 U18413 ( .A0(n8883), .A1(n8910), .S(n3318), .Z(N2861) );
  CMX2X1 U18414 ( .A0(mem_data1[800]), .A1(mem_data1[801]), .S(n4274), .Z(
        n8890) );
  CMXI2X1 U18415 ( .A0(n8890), .A1(n8884), .S(n4023), .Z(n8900) );
  CMX2X1 U18416 ( .A0(n8885), .A1(n8900), .S(n3796), .Z(n8913) );
  CMXI2X1 U18417 ( .A0(n8886), .A1(n8913), .S(n3318), .Z(N2862) );
  CMX2X1 U18418 ( .A0(mem_data1[801]), .A1(mem_data1[802]), .S(n4274), .Z(
        n8893) );
  CMXI2X1 U18419 ( .A0(n8893), .A1(n8887), .S(n4023), .Z(n8903) );
  CMX2X1 U18420 ( .A0(n8888), .A1(n8903), .S(n3797), .Z(n8916) );
  CMXI2X1 U18421 ( .A0(n8889), .A1(n8916), .S(n3318), .Z(N2863) );
  CMX2X1 U18422 ( .A0(mem_data1[802]), .A1(mem_data1[803]), .S(n4274), .Z(
        n8899) );
  CMXI2X1 U18423 ( .A0(n8899), .A1(n8890), .S(n4023), .Z(n8906) );
  CMX2X1 U18424 ( .A0(n8891), .A1(n8906), .S(n3805), .Z(n8919) );
  CMXI2X1 U18425 ( .A0(n8892), .A1(n8919), .S(n3318), .Z(N2864) );
  CMX2X1 U18426 ( .A0(mem_data1[803]), .A1(mem_data1[804]), .S(n4274), .Z(
        n8902) );
  CMXI2X1 U18427 ( .A0(n8902), .A1(n8893), .S(n4023), .Z(n8909) );
  CMX2X1 U18428 ( .A0(n8894), .A1(n8909), .S(n3806), .Z(n8922) );
  CMXI2X1 U18429 ( .A0(n8895), .A1(n8922), .S(n3318), .Z(N2865) );
  CMX2X1 U18430 ( .A0(mem_data1[92]), .A1(mem_data1[93]), .S(n4274), .Z(n8966)
         );
  CMXI2X1 U18431 ( .A0(n8966), .A1(n8896), .S(n4023), .Z(n9033) );
  CMX2X1 U18432 ( .A0(n8897), .A1(n9033), .S(n3807), .Z(n9167) );
  CMXI2X1 U18433 ( .A0(n8898), .A1(n9167), .S(n3318), .Z(N2154) );
  CMX2X1 U18434 ( .A0(mem_data1[804]), .A1(mem_data1[805]), .S(n4274), .Z(
        n8905) );
  CMXI2X1 U18435 ( .A0(n8905), .A1(n8899), .S(n4023), .Z(n8912) );
  CMX2X1 U18436 ( .A0(n8900), .A1(n8912), .S(n3808), .Z(n8925) );
  CMXI2X1 U18437 ( .A0(n8901), .A1(n8925), .S(n3318), .Z(N2866) );
  CMX2X1 U18438 ( .A0(mem_data1[805]), .A1(mem_data1[806]), .S(n4273), .Z(
        n8908) );
  CMXI2X1 U18439 ( .A0(n8908), .A1(n8902), .S(n4023), .Z(n8915) );
  CMX2X1 U18440 ( .A0(n8903), .A1(n8915), .S(n3809), .Z(n8928) );
  CMXI2X1 U18441 ( .A0(n8904), .A1(n8928), .S(n3318), .Z(N2867) );
  CMX2X1 U18442 ( .A0(mem_data1[806]), .A1(mem_data1[807]), .S(n4273), .Z(
        n8911) );
  CMXI2X1 U18443 ( .A0(n8911), .A1(n8905), .S(n4023), .Z(n8918) );
  CMX2X1 U18444 ( .A0(n8906), .A1(n8918), .S(n3810), .Z(n8938) );
  CMXI2X1 U18445 ( .A0(n8907), .A1(n8938), .S(n3318), .Z(N2868) );
  CMX2X1 U18446 ( .A0(mem_data1[807]), .A1(mem_data1[808]), .S(n4273), .Z(
        n8914) );
  CMXI2X1 U18447 ( .A0(n8914), .A1(n8908), .S(n4023), .Z(n8921) );
  CMX2X1 U18448 ( .A0(n8909), .A1(n8921), .S(n3811), .Z(n8941) );
  CMXI2X1 U18449 ( .A0(n8910), .A1(n8941), .S(n3318), .Z(N2869) );
  CMX2X1 U18450 ( .A0(mem_data1[808]), .A1(mem_data1[809]), .S(n4273), .Z(
        n8917) );
  CMXI2X1 U18451 ( .A0(n8917), .A1(n8911), .S(n4023), .Z(n8924) );
  CMX2X1 U18452 ( .A0(n8912), .A1(n8924), .S(n3812), .Z(n8944) );
  CMXI2X1 U18453 ( .A0(n8913), .A1(n8944), .S(n3317), .Z(N2870) );
  CMX2X1 U18454 ( .A0(mem_data1[809]), .A1(mem_data1[810]), .S(n4273), .Z(
        n8920) );
  CMXI2X1 U18455 ( .A0(n8920), .A1(n8914), .S(n4023), .Z(n8927) );
  CMX2X1 U18456 ( .A0(n8915), .A1(n8927), .S(n4361), .Z(n8947) );
  CMXI2X1 U18457 ( .A0(n8916), .A1(n8947), .S(n3317), .Z(N2871) );
  CMX2X1 U18458 ( .A0(mem_data1[810]), .A1(mem_data1[811]), .S(n4273), .Z(
        n8923) );
  CMXI2X1 U18459 ( .A0(n8923), .A1(n8917), .S(n4023), .Z(n8937) );
  CMX2X1 U18460 ( .A0(n8918), .A1(n8937), .S(n3771), .Z(n8950) );
  CMXI2X1 U18461 ( .A0(n8919), .A1(n8950), .S(n3317), .Z(N2872) );
  CMX2X1 U18462 ( .A0(mem_data1[811]), .A1(mem_data1[812]), .S(n4273), .Z(
        n8926) );
  CMXI2X1 U18463 ( .A0(n8926), .A1(n8920), .S(n4022), .Z(n8940) );
  CMX2X1 U18464 ( .A0(n8921), .A1(n8940), .S(n3773), .Z(n8953) );
  CMXI2X1 U18465 ( .A0(n8922), .A1(n8953), .S(n3317), .Z(N2873) );
  CMX2X1 U18466 ( .A0(mem_data1[812]), .A1(mem_data1[813]), .S(n4273), .Z(
        n8936) );
  CMXI2X1 U18467 ( .A0(n8936), .A1(n8923), .S(n4022), .Z(n8943) );
  CMX2X1 U18468 ( .A0(n8924), .A1(n8943), .S(n3772), .Z(n8956) );
  CMXI2X1 U18469 ( .A0(n8925), .A1(n8956), .S(n3317), .Z(N2874) );
  CMX2X1 U18470 ( .A0(mem_data1[813]), .A1(mem_data1[814]), .S(n4273), .Z(
        n8939) );
  CMXI2X1 U18471 ( .A0(n8939), .A1(n8926), .S(n4022), .Z(n8946) );
  CMX2X1 U18472 ( .A0(n8927), .A1(n8946), .S(n3774), .Z(n8959) );
  CMXI2X1 U18473 ( .A0(n8928), .A1(n8959), .S(n3317), .Z(N2875) );
  CMX2X1 U18474 ( .A0(mem_data1[93]), .A1(mem_data1[94]), .S(n4273), .Z(n8999)
         );
  CMXI2X1 U18475 ( .A0(n8999), .A1(n8929), .S(n4022), .Z(n9066) );
  CMX2X1 U18476 ( .A0(n8930), .A1(n9066), .S(n3775), .Z(n9201) );
  CMXI2X1 U18477 ( .A0(n8931), .A1(n9201), .S(n3320), .Z(N2155) );
  CMXI2X1 U18478 ( .A0(n4418), .A1(n8933), .S(n3781), .Z(n8935) );
  CMXI2X1 U18479 ( .A0(n8935), .A1(n8934), .S(n3320), .Z(N2083) );
  CMX2X1 U18480 ( .A0(mem_data1[814]), .A1(mem_data1[815]), .S(n4273), .Z(
        n8942) );
  CMXI2X1 U18481 ( .A0(n8942), .A1(n8936), .S(n4022), .Z(n8949) );
  CMX2X1 U18482 ( .A0(n8937), .A1(n8949), .S(n3776), .Z(n8962) );
  CMXI2X1 U18483 ( .A0(n8938), .A1(n8962), .S(n3320), .Z(N2876) );
  CMX2X1 U18484 ( .A0(mem_data1[815]), .A1(mem_data1[816]), .S(n4272), .Z(
        n8945) );
  CMXI2X1 U18485 ( .A0(n8945), .A1(n8939), .S(n4022), .Z(n8952) );
  CMX2X1 U18486 ( .A0(n8940), .A1(n8952), .S(n3777), .Z(n8965) );
  CMXI2X1 U18487 ( .A0(n8941), .A1(n8965), .S(n3320), .Z(N2877) );
  CMX2X1 U18488 ( .A0(mem_data1[816]), .A1(mem_data1[817]), .S(n4272), .Z(
        n8948) );
  CMXI2X1 U18489 ( .A0(n8948), .A1(n8942), .S(n4022), .Z(n8955) );
  CMX2X1 U18490 ( .A0(n8943), .A1(n8955), .S(n3790), .Z(n8971) );
  CMXI2X1 U18491 ( .A0(n8944), .A1(n8971), .S(n3320), .Z(N2878) );
  CMX2X1 U18492 ( .A0(mem_data1[817]), .A1(mem_data1[818]), .S(n4272), .Z(
        n8951) );
  CMXI2X1 U18493 ( .A0(n8951), .A1(n8945), .S(n4022), .Z(n8958) );
  CMX2X1 U18494 ( .A0(n8946), .A1(n8958), .S(n3796), .Z(n8974) );
  CMXI2X1 U18495 ( .A0(n8947), .A1(n8974), .S(n3320), .Z(N2879) );
  CMX2X1 U18496 ( .A0(mem_data1[818]), .A1(mem_data1[819]), .S(n4272), .Z(
        n8954) );
  CMXI2X1 U18497 ( .A0(n8954), .A1(n8948), .S(n4022), .Z(n8961) );
  CMX2X1 U18498 ( .A0(n8949), .A1(n8961), .S(n3772), .Z(n8977) );
  CMXI2X1 U18499 ( .A0(n8950), .A1(n8977), .S(n3320), .Z(N2880) );
  CMX2X1 U18500 ( .A0(mem_data1[819]), .A1(mem_data1[820]), .S(n4272), .Z(
        n8957) );
  CMXI2X1 U18501 ( .A0(n8957), .A1(n8951), .S(n4022), .Z(n8964) );
  CMX2X1 U18502 ( .A0(n8952), .A1(n8964), .S(n3773), .Z(n8980) );
  CMXI2X1 U18503 ( .A0(n8953), .A1(n8980), .S(n3320), .Z(N2881) );
  CMX2X1 U18504 ( .A0(mem_data1[820]), .A1(mem_data1[821]), .S(n4272), .Z(
        n8960) );
  CMXI2X1 U18505 ( .A0(n8960), .A1(n8954), .S(n4022), .Z(n8970) );
  CMX2X1 U18506 ( .A0(n8955), .A1(n8970), .S(n3774), .Z(n8983) );
  CMXI2X1 U18507 ( .A0(n8956), .A1(n8983), .S(n3319), .Z(N2882) );
  CMX2X1 U18508 ( .A0(mem_data1[821]), .A1(mem_data1[822]), .S(n4272), .Z(
        n8963) );
  CMXI2X1 U18509 ( .A0(n8963), .A1(n8957), .S(n4022), .Z(n8973) );
  CMX2X1 U18510 ( .A0(n8958), .A1(n8973), .S(n3775), .Z(n8986) );
  CMXI2X1 U18511 ( .A0(n8959), .A1(n8986), .S(n3319), .Z(N2883) );
  CMX2X1 U18512 ( .A0(mem_data1[822]), .A1(mem_data1[823]), .S(n4272), .Z(
        n8969) );
  CMXI2X1 U18513 ( .A0(n8969), .A1(n8960), .S(n4022), .Z(n8976) );
  CMX2X1 U18514 ( .A0(n8961), .A1(n8976), .S(n3776), .Z(n8989) );
  CMXI2X1 U18515 ( .A0(n8962), .A1(n8989), .S(n3319), .Z(N2884) );
  CMX2X1 U18516 ( .A0(mem_data1[823]), .A1(mem_data1[824]), .S(n4272), .Z(
        n8972) );
  CMXI2X1 U18517 ( .A0(n8972), .A1(n8963), .S(n4022), .Z(n8979) );
  CMX2X1 U18518 ( .A0(n8964), .A1(n8979), .S(n3777), .Z(n8992) );
  CMXI2X1 U18519 ( .A0(n8965), .A1(n8992), .S(n3319), .Z(N2885) );
  CMX2X1 U18520 ( .A0(mem_data1[94]), .A1(mem_data1[95]), .S(n4272), .Z(n9032)
         );
  CMXI2X1 U18521 ( .A0(n9032), .A1(n8966), .S(n4022), .Z(n9099) );
  CMX2X1 U18522 ( .A0(n8967), .A1(n9099), .S(n3790), .Z(n9234) );
  CMXI2X1 U18523 ( .A0(n8968), .A1(n9234), .S(n3319), .Z(N2156) );
  CMX2X1 U18524 ( .A0(mem_data1[824]), .A1(mem_data1[825]), .S(n4272), .Z(
        n8975) );
  CMXI2X1 U18525 ( .A0(n8975), .A1(n8969), .S(n4022), .Z(n8982) );
  CMX2X1 U18526 ( .A0(n8970), .A1(n8982), .S(n3791), .Z(n8995) );
  CMXI2X1 U18527 ( .A0(n8971), .A1(n8995), .S(n3319), .Z(N2886) );
  CMX2X1 U18528 ( .A0(mem_data1[825]), .A1(mem_data1[826]), .S(n4271), .Z(
        n8978) );
  CMXI2X1 U18529 ( .A0(n8978), .A1(n8972), .S(n4021), .Z(n8985) );
  CMX2X1 U18530 ( .A0(n8973), .A1(n8985), .S(n3792), .Z(n8998) );
  CMXI2X1 U18531 ( .A0(n8974), .A1(n8998), .S(n3319), .Z(N2887) );
  CMX2X1 U18532 ( .A0(mem_data1[826]), .A1(mem_data1[827]), .S(n4271), .Z(
        n8981) );
  CMXI2X1 U18533 ( .A0(n8981), .A1(n8975), .S(n4021), .Z(n8988) );
  CMX2X1 U18534 ( .A0(n8976), .A1(n8988), .S(n3793), .Z(n9004) );
  CMXI2X1 U18535 ( .A0(n8977), .A1(n9004), .S(n3319), .Z(N2888) );
  CMX2X1 U18536 ( .A0(mem_data1[827]), .A1(mem_data1[828]), .S(n4271), .Z(
        n8984) );
  CMXI2X1 U18537 ( .A0(n8984), .A1(n8978), .S(n4021), .Z(n8991) );
  CMX2X1 U18538 ( .A0(n8979), .A1(n8991), .S(n3794), .Z(n9007) );
  CMXI2X1 U18539 ( .A0(n8980), .A1(n9007), .S(n3319), .Z(N2889) );
  CMX2X1 U18540 ( .A0(mem_data1[828]), .A1(mem_data1[829]), .S(n4271), .Z(
        n8987) );
  CMXI2X1 U18541 ( .A0(n8987), .A1(n8981), .S(n4021), .Z(n8994) );
  CMX2X1 U18542 ( .A0(n8982), .A1(n8994), .S(n3795), .Z(n9010) );
  CMXI2X1 U18543 ( .A0(n8983), .A1(n9010), .S(n3319), .Z(N2890) );
  CMX2X1 U18544 ( .A0(mem_data1[829]), .A1(mem_data1[830]), .S(n4271), .Z(
        n8990) );
  CMXI2X1 U18545 ( .A0(n8990), .A1(n8984), .S(n4021), .Z(n8997) );
  CMX2X1 U18546 ( .A0(n8985), .A1(n8997), .S(n3796), .Z(n9013) );
  CMXI2X1 U18547 ( .A0(n8986), .A1(n9013), .S(n3322), .Z(N2891) );
  CMX2X1 U18548 ( .A0(mem_data1[830]), .A1(mem_data1[831]), .S(n4271), .Z(
        n8993) );
  CMXI2X1 U18549 ( .A0(n8993), .A1(n8987), .S(n4021), .Z(n9003) );
  CMX2X1 U18550 ( .A0(n8988), .A1(n9003), .S(n3797), .Z(n9016) );
  CMXI2X1 U18551 ( .A0(n8989), .A1(n9016), .S(n3322), .Z(N2892) );
  CMX2X1 U18552 ( .A0(mem_data1[831]), .A1(mem_data1[832]), .S(n4271), .Z(
        n8996) );
  CMXI2X1 U18553 ( .A0(n8996), .A1(n8990), .S(n4021), .Z(n9006) );
  CMX2X1 U18554 ( .A0(n8991), .A1(n9006), .S(n3805), .Z(n9019) );
  CMXI2X1 U18555 ( .A0(n8992), .A1(n9019), .S(n3322), .Z(N2893) );
  CMX2X1 U18556 ( .A0(mem_data1[832]), .A1(mem_data1[833]), .S(n4271), .Z(
        n9002) );
  CMXI2X1 U18557 ( .A0(n9002), .A1(n8993), .S(n4021), .Z(n9009) );
  CMX2X1 U18558 ( .A0(n8994), .A1(n9009), .S(n3806), .Z(n9022) );
  CMXI2X1 U18559 ( .A0(n8995), .A1(n9022), .S(n3322), .Z(N2894) );
  CMX2X1 U18560 ( .A0(mem_data1[833]), .A1(mem_data1[834]), .S(n4271), .Z(
        n9005) );
  CMXI2X1 U18561 ( .A0(n9005), .A1(n8996), .S(n4021), .Z(n9012) );
  CMX2X1 U18562 ( .A0(n8997), .A1(n9012), .S(n3774), .Z(n9025) );
  CMXI2X1 U18563 ( .A0(n8998), .A1(n9025), .S(n3321), .Z(N2895) );
  CMX2X1 U18564 ( .A0(mem_data1[95]), .A1(mem_data1[96]), .S(n4271), .Z(n9065)
         );
  CMXI2X1 U18565 ( .A0(n9065), .A1(n8999), .S(n4021), .Z(n9132) );
  CMX2X1 U18566 ( .A0(n9000), .A1(n9132), .S(n3773), .Z(n9267) );
  CMXI2X1 U18567 ( .A0(n9001), .A1(n9267), .S(n3321), .Z(N2157) );
  CMX2X1 U18568 ( .A0(mem_data1[834]), .A1(mem_data1[835]), .S(n4271), .Z(
        n9008) );
  CMXI2X1 U18569 ( .A0(n9008), .A1(n9002), .S(n4021), .Z(n9015) );
  CMX2X1 U18570 ( .A0(n9003), .A1(n9015), .S(n3791), .Z(n9028) );
  CMXI2X1 U18571 ( .A0(n9004), .A1(n9028), .S(n3321), .Z(N2896) );
  CMX2X1 U18572 ( .A0(mem_data1[835]), .A1(mem_data1[836]), .S(n4270), .Z(
        n9011) );
  CMXI2X1 U18573 ( .A0(n9011), .A1(n9005), .S(n4021), .Z(n9018) );
  CMX2X1 U18574 ( .A0(n9006), .A1(n9018), .S(n3792), .Z(n9031) );
  CMXI2X1 U18575 ( .A0(n9007), .A1(n9031), .S(n3321), .Z(N2897) );
  CMX2X1 U18576 ( .A0(mem_data1[836]), .A1(mem_data1[837]), .S(n4270), .Z(
        n9014) );
  CMXI2X1 U18577 ( .A0(n9014), .A1(n9008), .S(n4021), .Z(n9021) );
  CMX2X1 U18578 ( .A0(n9009), .A1(n9021), .S(n3793), .Z(n9037) );
  CMXI2X1 U18579 ( .A0(n9010), .A1(n9037), .S(n3321), .Z(N2898) );
  CMX2X1 U18580 ( .A0(mem_data1[837]), .A1(mem_data1[838]), .S(n4270), .Z(
        n9017) );
  CMXI2X1 U18581 ( .A0(n9017), .A1(n9011), .S(n4021), .Z(n9024) );
  CMX2X1 U18582 ( .A0(n9012), .A1(n9024), .S(n3794), .Z(n9040) );
  CMXI2X1 U18583 ( .A0(n9013), .A1(n9040), .S(n3321), .Z(N2899) );
  CMX2X1 U18584 ( .A0(mem_data1[838]), .A1(mem_data1[839]), .S(n4270), .Z(
        n9020) );
  CMXI2X1 U18585 ( .A0(n9020), .A1(n9014), .S(n4021), .Z(n9027) );
  CMX2X1 U18586 ( .A0(n9015), .A1(n9027), .S(n3795), .Z(n9043) );
  CMXI2X1 U18587 ( .A0(n9016), .A1(n9043), .S(n3321), .Z(N2900) );
  CMX2X1 U18588 ( .A0(mem_data1[839]), .A1(mem_data1[840]), .S(n4270), .Z(
        n9023) );
  CMXI2X1 U18589 ( .A0(n9023), .A1(n9017), .S(n4021), .Z(n9030) );
  CMX2X1 U18590 ( .A0(n9018), .A1(n9030), .S(n3797), .Z(n9046) );
  CMXI2X1 U18591 ( .A0(n9019), .A1(n9046), .S(n3321), .Z(N2901) );
  CMX2X1 U18592 ( .A0(mem_data1[840]), .A1(mem_data1[841]), .S(n4270), .Z(
        n9026) );
  CMXI2X1 U18593 ( .A0(n9026), .A1(n9020), .S(n4020), .Z(n9036) );
  CMX2X1 U18594 ( .A0(n9021), .A1(n9036), .S(n3807), .Z(n9049) );
  CMXI2X1 U18595 ( .A0(n9022), .A1(n9049), .S(n3321), .Z(N2902) );
  CMX2X1 U18596 ( .A0(mem_data1[841]), .A1(mem_data1[842]), .S(n4270), .Z(
        n9029) );
  CMXI2X1 U18597 ( .A0(n9029), .A1(n9023), .S(n4020), .Z(n9039) );
  CMX2X1 U18598 ( .A0(n9024), .A1(n9039), .S(n3808), .Z(n9052) );
  CMXI2X1 U18599 ( .A0(n9025), .A1(n9052), .S(n3321), .Z(N2903) );
  CMX2X1 U18600 ( .A0(mem_data1[842]), .A1(mem_data1[843]), .S(n4270), .Z(
        n9035) );
  CMXI2X1 U18601 ( .A0(n9035), .A1(n9026), .S(n4020), .Z(n9042) );
  CMX2X1 U18602 ( .A0(n9027), .A1(n9042), .S(n3809), .Z(n9055) );
  CMXI2X1 U18603 ( .A0(n9028), .A1(n9055), .S(n3321), .Z(N2904) );
  CMX2X1 U18604 ( .A0(mem_data1[843]), .A1(mem_data1[844]), .S(n4278), .Z(
        n9038) );
  CMXI2X1 U18605 ( .A0(n9038), .A1(n9029), .S(n4020), .Z(n9045) );
  CMX2X1 U18606 ( .A0(n9030), .A1(n9045), .S(n3810), .Z(n9058) );
  CMXI2X1 U18607 ( .A0(n9031), .A1(n9058), .S(n3320), .Z(N2905) );
  CMX2X1 U18608 ( .A0(mem_data1[96]), .A1(mem_data1[97]), .S(n4270), .Z(n9098)
         );
  CMXI2X1 U18609 ( .A0(n9098), .A1(n9032), .S(n4020), .Z(n9166) );
  CMX2X1 U18610 ( .A0(n9033), .A1(n9166), .S(n3811), .Z(n9302) );
  CMXI2X1 U18611 ( .A0(n9034), .A1(n9302), .S(n3320), .Z(N2158) );
  CMX2X1 U18612 ( .A0(mem_data1[844]), .A1(mem_data1[845]), .S(n4270), .Z(
        n9041) );
  CMXI2X1 U18613 ( .A0(n9041), .A1(n9035), .S(n4020), .Z(n9048) );
  CMX2X1 U18614 ( .A0(n9036), .A1(n9048), .S(n3812), .Z(n9061) );
  CMXI2X1 U18615 ( .A0(n9037), .A1(n9061), .S(n3320), .Z(N2906) );
  CMX2X1 U18616 ( .A0(mem_data1[845]), .A1(mem_data1[846]), .S(n4269), .Z(
        n9044) );
  CMXI2X1 U18617 ( .A0(n9044), .A1(n9038), .S(n4020), .Z(n9051) );
  CMX2X1 U18618 ( .A0(n9039), .A1(n9051), .S(n4358), .Z(n9064) );
  CMXI2X1 U18619 ( .A0(n9040), .A1(n9064), .S(n3323), .Z(N2907) );
  CMX2X1 U18620 ( .A0(mem_data1[846]), .A1(mem_data1[847]), .S(n4269), .Z(
        n9047) );
  CMXI2X1 U18621 ( .A0(n9047), .A1(n9041), .S(n4020), .Z(n9054) );
  CMX2X1 U18622 ( .A0(n9042), .A1(n9054), .S(n3771), .Z(n9070) );
  CMXI2X1 U18623 ( .A0(n9043), .A1(n9070), .S(n3323), .Z(N2908) );
  CMX2X1 U18624 ( .A0(mem_data1[847]), .A1(mem_data1[848]), .S(n4269), .Z(
        n9050) );
  CMXI2X1 U18625 ( .A0(n9050), .A1(n9044), .S(n4020), .Z(n9057) );
  CMX2X1 U18626 ( .A0(n9045), .A1(n9057), .S(n3772), .Z(n9073) );
  CMXI2X1 U18627 ( .A0(n9046), .A1(n9073), .S(n3323), .Z(N2909) );
  CMX2X1 U18628 ( .A0(mem_data1[848]), .A1(mem_data1[849]), .S(n4269), .Z(
        n9053) );
  CMXI2X1 U18629 ( .A0(n9053), .A1(n9047), .S(n4020), .Z(n9060) );
  CMX2X1 U18630 ( .A0(n9048), .A1(n9060), .S(n3773), .Z(n9076) );
  CMXI2X1 U18631 ( .A0(n9049), .A1(n9076), .S(n3323), .Z(N2910) );
  CMX2X1 U18632 ( .A0(mem_data1[849]), .A1(mem_data1[850]), .S(n4269), .Z(
        n9056) );
  CMXI2X1 U18633 ( .A0(n9056), .A1(n9050), .S(n4020), .Z(n9063) );
  CMX2X1 U18634 ( .A0(n9051), .A1(n9063), .S(n3774), .Z(n9079) );
  CMXI2X1 U18635 ( .A0(n9052), .A1(n9079), .S(n3323), .Z(N2911) );
  CMX2X1 U18636 ( .A0(mem_data1[850]), .A1(mem_data1[851]), .S(n4269), .Z(
        n9059) );
  CMXI2X1 U18637 ( .A0(n9059), .A1(n9053), .S(n4020), .Z(n9069) );
  CMX2X1 U18638 ( .A0(n9054), .A1(n9069), .S(n3775), .Z(n9082) );
  CMXI2X1 U18639 ( .A0(n9055), .A1(n9082), .S(n3323), .Z(N2912) );
  CMX2X1 U18640 ( .A0(mem_data1[851]), .A1(mem_data1[852]), .S(n4269), .Z(
        n9062) );
  CMXI2X1 U18641 ( .A0(n9062), .A1(n9056), .S(n4020), .Z(n9072) );
  CMX2X1 U18642 ( .A0(n9057), .A1(n9072), .S(n3776), .Z(n9085) );
  CMXI2X1 U18643 ( .A0(n9058), .A1(n9085), .S(n3323), .Z(N2913) );
  CMX2X1 U18644 ( .A0(mem_data1[852]), .A1(mem_data1[853]), .S(n4269), .Z(
        n9068) );
  CMXI2X1 U18645 ( .A0(n9068), .A1(n9059), .S(n4020), .Z(n9075) );
  CMX2X1 U18646 ( .A0(n9060), .A1(n9075), .S(n3777), .Z(n9088) );
  CMXI2X1 U18647 ( .A0(n9061), .A1(n9088), .S(n3323), .Z(N2914) );
  CMX2X1 U18648 ( .A0(mem_data1[853]), .A1(mem_data1[854]), .S(n4269), .Z(
        n9071) );
  CMXI2X1 U18649 ( .A0(n9071), .A1(n9062), .S(n4020), .Z(n9078) );
  CMX2X1 U18650 ( .A0(n9063), .A1(n9078), .S(n3790), .Z(n9091) );
  CMXI2X1 U18651 ( .A0(n9064), .A1(n9091), .S(n3323), .Z(N2915) );
  CMX2X1 U18652 ( .A0(mem_data1[97]), .A1(mem_data1[98]), .S(n4269), .Z(n9131)
         );
  CMXI2X1 U18653 ( .A0(n9131), .A1(n9065), .S(n4020), .Z(n9200) );
  CMX2X1 U18654 ( .A0(n9066), .A1(n9200), .S(n3791), .Z(n9335) );
  CMXI2X1 U18655 ( .A0(n9067), .A1(n9335), .S(n3323), .Z(N2159) );
  CMX2X1 U18656 ( .A0(mem_data1[854]), .A1(mem_data1[855]), .S(n4269), .Z(
        n9074) );
  CMXI2X1 U18657 ( .A0(n9074), .A1(n9068), .S(n4019), .Z(n9081) );
  CMX2X1 U18658 ( .A0(n9069), .A1(n9081), .S(n3775), .Z(n9094) );
  CMXI2X1 U18659 ( .A0(n9070), .A1(n9094), .S(n3323), .Z(N2916) );
  CMX2X1 U18660 ( .A0(mem_data1[855]), .A1(mem_data1[856]), .S(n4268), .Z(
        n9077) );
  CMXI2X1 U18661 ( .A0(n9077), .A1(n9071), .S(n4019), .Z(n9084) );
  CMX2X1 U18662 ( .A0(n9072), .A1(n9084), .S(n3774), .Z(n9097) );
  CMXI2X1 U18663 ( .A0(n9073), .A1(n9097), .S(n3322), .Z(N2917) );
  CMX2X1 U18664 ( .A0(mem_data1[856]), .A1(mem_data1[857]), .S(n4268), .Z(
        n9080) );
  CMXI2X1 U18665 ( .A0(n9080), .A1(n9074), .S(n4019), .Z(n9087) );
  CMX2X1 U18666 ( .A0(n9075), .A1(n9087), .S(n3797), .Z(n9103) );
  CMXI2X1 U18667 ( .A0(n9076), .A1(n9103), .S(n3322), .Z(N2918) );
  CMX2X1 U18668 ( .A0(mem_data1[857]), .A1(mem_data1[858]), .S(n4268), .Z(
        n9083) );
  CMXI2X1 U18669 ( .A0(n9083), .A1(n9077), .S(n4019), .Z(n9090) );
  CMX2X1 U18670 ( .A0(n9078), .A1(n9090), .S(n3805), .Z(n9106) );
  CMXI2X1 U18671 ( .A0(n9079), .A1(n9106), .S(n3322), .Z(N2919) );
  CMX2X1 U18672 ( .A0(mem_data1[858]), .A1(mem_data1[859]), .S(n4268), .Z(
        n9086) );
  CMXI2X1 U18673 ( .A0(n9086), .A1(n9080), .S(n4019), .Z(n9093) );
  CMX2X1 U18674 ( .A0(n9081), .A1(n9093), .S(n3806), .Z(n9109) );
  CMXI2X1 U18675 ( .A0(n9082), .A1(n9109), .S(n3322), .Z(N2920) );
  CMX2X1 U18676 ( .A0(mem_data1[859]), .A1(mem_data1[860]), .S(n4268), .Z(
        n9089) );
  CMXI2X1 U18677 ( .A0(n9089), .A1(n9083), .S(n4019), .Z(n9096) );
  CMX2X1 U18678 ( .A0(n9084), .A1(n9096), .S(n3808), .Z(n9112) );
  CMXI2X1 U18679 ( .A0(n9085), .A1(n9112), .S(n3322), .Z(N2921) );
  CMX2X1 U18680 ( .A0(mem_data1[860]), .A1(mem_data1[861]), .S(n4268), .Z(
        n9092) );
  CMXI2X1 U18681 ( .A0(n9092), .A1(n9086), .S(n4019), .Z(n9102) );
  CMX2X1 U18682 ( .A0(n9087), .A1(n9102), .S(n3809), .Z(n9115) );
  CMXI2X1 U18683 ( .A0(n9088), .A1(n9115), .S(n3322), .Z(N2922) );
  CMX2X1 U18684 ( .A0(mem_data1[861]), .A1(mem_data1[862]), .S(n4268), .Z(
        n9095) );
  CMXI2X1 U18685 ( .A0(n9095), .A1(n9089), .S(n4019), .Z(n9105) );
  CMX2X1 U18686 ( .A0(n9090), .A1(n9105), .S(n3812), .Z(n9118) );
  CMXI2X1 U18687 ( .A0(n9091), .A1(n9118), .S(n3322), .Z(N2923) );
  CMX2X1 U18688 ( .A0(mem_data1[862]), .A1(mem_data1[863]), .S(n4268), .Z(
        n9101) );
  CMXI2X1 U18689 ( .A0(n9101), .A1(n9092), .S(n4019), .Z(n9108) );
  CMX2X1 U18690 ( .A0(n9093), .A1(n9108), .S(n3772), .Z(n9121) );
  CMXI2X1 U18691 ( .A0(n9094), .A1(n9121), .S(n3325), .Z(N2924) );
  CMX2X1 U18692 ( .A0(mem_data1[863]), .A1(mem_data1[864]), .S(n4268), .Z(
        n9104) );
  CMXI2X1 U18693 ( .A0(n9104), .A1(n9095), .S(n4019), .Z(n9111) );
  CMX2X1 U18694 ( .A0(n9096), .A1(n9111), .S(n3773), .Z(n9124) );
  CMXI2X1 U18695 ( .A0(n9097), .A1(n9124), .S(n3325), .Z(N2925) );
  CMX2X1 U18696 ( .A0(mem_data1[98]), .A1(mem_data1[99]), .S(n4268), .Z(n9164)
         );
  CMXI2X1 U18697 ( .A0(n9164), .A1(n9098), .S(n4019), .Z(n9233) );
  CMX2X1 U18698 ( .A0(n9099), .A1(n9233), .S(n3774), .Z(n9367) );
  CMXI2X1 U18699 ( .A0(n9100), .A1(n9367), .S(n3325), .Z(N2160) );
  CMX2X1 U18700 ( .A0(mem_data1[864]), .A1(mem_data1[865]), .S(n4268), .Z(
        n9107) );
  CMXI2X1 U18701 ( .A0(n9107), .A1(n9101), .S(n4019), .Z(n9114) );
  CMX2X1 U18702 ( .A0(n9102), .A1(n9114), .S(n3775), .Z(n9127) );
  CMXI2X1 U18703 ( .A0(n9103), .A1(n9127), .S(n3325), .Z(N2926) );
  CMX2X1 U18704 ( .A0(mem_data1[865]), .A1(mem_data1[866]), .S(n4267), .Z(
        n9110) );
  CMXI2X1 U18705 ( .A0(n9110), .A1(n9104), .S(n4019), .Z(n9117) );
  CMX2X1 U18706 ( .A0(n9105), .A1(n9117), .S(n3776), .Z(n9130) );
  CMXI2X1 U18707 ( .A0(n9106), .A1(n9130), .S(n3325), .Z(N2927) );
  CMX2X1 U18708 ( .A0(mem_data1[866]), .A1(mem_data1[867]), .S(n4267), .Z(
        n9113) );
  CMXI2X1 U18709 ( .A0(n9113), .A1(n9107), .S(n4019), .Z(n9120) );
  CMX2X1 U18710 ( .A0(n9108), .A1(n9120), .S(n3777), .Z(n9136) );
  CMXI2X1 U18711 ( .A0(n9109), .A1(n9136), .S(n3325), .Z(N2928) );
  CMX2X1 U18712 ( .A0(mem_data1[867]), .A1(mem_data1[868]), .S(n4267), .Z(
        n9116) );
  CMXI2X1 U18713 ( .A0(n9116), .A1(n9110), .S(n4019), .Z(n9123) );
  CMX2X1 U18714 ( .A0(n9111), .A1(n9123), .S(n3790), .Z(n9139) );
  CMXI2X1 U18715 ( .A0(n9112), .A1(n9139), .S(n3325), .Z(N2929) );
  CMX2X1 U18716 ( .A0(mem_data1[868]), .A1(mem_data1[869]), .S(n4267), .Z(
        n9119) );
  CMXI2X1 U18717 ( .A0(n9119), .A1(n9113), .S(n4019), .Z(n9126) );
  CMX2X1 U18718 ( .A0(n9114), .A1(n9126), .S(n3791), .Z(n9142) );
  CMXI2X1 U18719 ( .A0(n9115), .A1(n9142), .S(n3324), .Z(N2930) );
  CMX2X1 U18720 ( .A0(mem_data1[869]), .A1(mem_data1[870]), .S(n4267), .Z(
        n9122) );
  CMXI2X1 U18721 ( .A0(n9122), .A1(n9116), .S(n4018), .Z(n9129) );
  CMX2X1 U18722 ( .A0(n9117), .A1(n9129), .S(n3792), .Z(n9145) );
  CMXI2X1 U18723 ( .A0(n9118), .A1(n9145), .S(n3324), .Z(N2931) );
  CMX2X1 U18724 ( .A0(mem_data1[870]), .A1(mem_data1[871]), .S(n4267), .Z(
        n9125) );
  CMXI2X1 U18725 ( .A0(n9125), .A1(n9119), .S(n4018), .Z(n9135) );
  CMX2X1 U18726 ( .A0(n9120), .A1(n9135), .S(n3793), .Z(n9148) );
  CMXI2X1 U18727 ( .A0(n9121), .A1(n9148), .S(n3324), .Z(N2932) );
  CMX2X1 U18728 ( .A0(mem_data1[871]), .A1(mem_data1[872]), .S(n4267), .Z(
        n9128) );
  CMXI2X1 U18729 ( .A0(n9128), .A1(n9122), .S(n4018), .Z(n9138) );
  CMX2X1 U18730 ( .A0(n9123), .A1(n9138), .S(n3794), .Z(n9151) );
  CMXI2X1 U18731 ( .A0(n9124), .A1(n9151), .S(n3324), .Z(N2933) );
  CMX2X1 U18732 ( .A0(mem_data1[872]), .A1(mem_data1[873]), .S(n4267), .Z(
        n9134) );
  CMXI2X1 U18733 ( .A0(n9134), .A1(n9125), .S(n4018), .Z(n9141) );
  CMX2X1 U18734 ( .A0(n9126), .A1(n9141), .S(n3795), .Z(n9154) );
  CMXI2X1 U18735 ( .A0(n9127), .A1(n9154), .S(n3324), .Z(N2934) );
  CMX2X1 U18736 ( .A0(mem_data1[873]), .A1(mem_data1[874]), .S(n4267), .Z(
        n9137) );
  CMXI2X1 U18737 ( .A0(n9137), .A1(n9128), .S(n4018), .Z(n9144) );
  CMX2X1 U18738 ( .A0(n9129), .A1(n9144), .S(n3796), .Z(n9157) );
  CMXI2X1 U18739 ( .A0(n9130), .A1(n9157), .S(n3324), .Z(N2935) );
  CMX2X1 U18740 ( .A0(mem_data1[99]), .A1(mem_data1[100]), .S(n4267), .Z(n9198) );
  CMXI2X1 U18741 ( .A0(n9198), .A1(n9131), .S(n4018), .Z(n9266) );
  CMX2X1 U18742 ( .A0(n9132), .A1(n9266), .S(n3797), .Z(n9399) );
  CMXI2X1 U18743 ( .A0(n9133), .A1(n9399), .S(n3324), .Z(N2161) );
  CMX2X1 U18744 ( .A0(mem_data1[874]), .A1(mem_data1[875]), .S(n4267), .Z(
        n9140) );
  CMXI2X1 U18745 ( .A0(n9140), .A1(n9134), .S(n4018), .Z(n9147) );
  CMX2X1 U18746 ( .A0(n9135), .A1(n9147), .S(n3805), .Z(n9160) );
  CMXI2X1 U18747 ( .A0(n9136), .A1(n9160), .S(n3324), .Z(N2936) );
  CMX2X1 U18748 ( .A0(mem_data1[875]), .A1(mem_data1[876]), .S(n4266), .Z(
        n9143) );
  CMXI2X1 U18749 ( .A0(n9143), .A1(n9137), .S(n4018), .Z(n9150) );
  CMX2X1 U18750 ( .A0(n9138), .A1(n9150), .S(n3806), .Z(n9163) );
  CMXI2X1 U18751 ( .A0(n9139), .A1(n9163), .S(n3324), .Z(N2937) );
  CMX2X1 U18752 ( .A0(mem_data1[876]), .A1(mem_data1[877]), .S(n4266), .Z(
        n9146) );
  CMXI2X1 U18753 ( .A0(n9146), .A1(n9140), .S(n4018), .Z(n9153) );
  CMX2X1 U18754 ( .A0(n9141), .A1(n9153), .S(n3772), .Z(n9170) );
  CMXI2X1 U18755 ( .A0(n9142), .A1(n9170), .S(n3324), .Z(N2938) );
  CMX2X1 U18756 ( .A0(mem_data1[877]), .A1(mem_data1[878]), .S(n4266), .Z(
        n9149) );
  CMXI2X1 U18757 ( .A0(n9149), .A1(n9143), .S(n4018), .Z(n9156) );
  CMX2X1 U18758 ( .A0(n9144), .A1(n9156), .S(n3792), .Z(n9173) );
  CMXI2X1 U18759 ( .A0(n9145), .A1(n9173), .S(n3327), .Z(N2939) );
  CMX2X1 U18760 ( .A0(mem_data1[878]), .A1(mem_data1[879]), .S(n4266), .Z(
        n9152) );
  CMXI2X1 U18761 ( .A0(n9152), .A1(n9146), .S(n4018), .Z(n9159) );
  CMX2X1 U18762 ( .A0(n9147), .A1(n9159), .S(n3810), .Z(n9176) );
  CMXI2X1 U18763 ( .A0(n9148), .A1(n9176), .S(n3327), .Z(N2940) );
  CMX2X1 U18764 ( .A0(mem_data1[879]), .A1(mem_data1[880]), .S(n4266), .Z(
        n9155) );
  CMXI2X1 U18765 ( .A0(n9155), .A1(n9149), .S(n4018), .Z(n9162) );
  CMX2X1 U18766 ( .A0(n9150), .A1(n9162), .S(n3777), .Z(n9179) );
  CMXI2X1 U18767 ( .A0(n9151), .A1(n9179), .S(n3327), .Z(N2941) );
  CMX2X1 U18768 ( .A0(mem_data1[880]), .A1(mem_data1[881]), .S(n4266), .Z(
        n9158) );
  CMXI2X1 U18769 ( .A0(n9158), .A1(n9152), .S(n4018), .Z(n9169) );
  CMX2X1 U18770 ( .A0(n9153), .A1(n9169), .S(n3791), .Z(n9182) );
  CMXI2X1 U18771 ( .A0(n9154), .A1(n9182), .S(n3327), .Z(N2942) );
  CMX2X1 U18772 ( .A0(mem_data1[881]), .A1(mem_data1[882]), .S(n4266), .Z(
        n9161) );
  CMXI2X1 U18773 ( .A0(n9161), .A1(n9155), .S(n4018), .Z(n9172) );
  CMX2X1 U18774 ( .A0(n9156), .A1(n9172), .S(n3807), .Z(n9185) );
  CMXI2X1 U18775 ( .A0(n9157), .A1(n9185), .S(n3326), .Z(N2943) );
  CMX2X1 U18776 ( .A0(mem_data1[882]), .A1(mem_data1[883]), .S(n4266), .Z(
        n9168) );
  CMXI2X1 U18777 ( .A0(n9168), .A1(n9158), .S(n4018), .Z(n9175) );
  CMX2X1 U18778 ( .A0(n9159), .A1(n9175), .S(n3808), .Z(n9188) );
  CMXI2X1 U18779 ( .A0(n9160), .A1(n9188), .S(n3326), .Z(N2944) );
  CMX2X1 U18780 ( .A0(mem_data1[883]), .A1(mem_data1[884]), .S(n4266), .Z(
        n9171) );
  CMXI2X1 U18781 ( .A0(n9171), .A1(n9161), .S(n4018), .Z(n9178) );
  CMX2X1 U18782 ( .A0(n9162), .A1(n9178), .S(n3809), .Z(n9191) );
  CMXI2X1 U18783 ( .A0(n9163), .A1(n9191), .S(n3326), .Z(N2945) );
  CMXI2X1 U18784 ( .A0(n9165), .A1(n9164), .S(n4017), .Z(n9301) );
  CMX2X1 U18785 ( .A0(n9166), .A1(n9301), .S(n3810), .Z(n9431) );
  CMXI2X1 U18786 ( .A0(n9167), .A1(n9431), .S(n3326), .Z(N2162) );
  CMX2X1 U18787 ( .A0(mem_data1[884]), .A1(mem_data1[885]), .S(n4266), .Z(
        n9174) );
  CMXI2X1 U18788 ( .A0(n9174), .A1(n9168), .S(n4017), .Z(n9181) );
  CMX2X1 U18789 ( .A0(n9169), .A1(n9181), .S(n3811), .Z(n9194) );
  CMXI2X1 U18790 ( .A0(n9170), .A1(n9194), .S(n3326), .Z(N2946) );
  CMX2X1 U18791 ( .A0(mem_data1[885]), .A1(mem_data1[886]), .S(n4266), .Z(
        n9177) );
  CMXI2X1 U18792 ( .A0(n9177), .A1(n9171), .S(n4017), .Z(n9184) );
  CMX2X1 U18793 ( .A0(n9172), .A1(n9184), .S(n3812), .Z(n9197) );
  CMXI2X1 U18794 ( .A0(n9173), .A1(n9197), .S(n3326), .Z(N2947) );
  CMX2X1 U18795 ( .A0(mem_data1[886]), .A1(mem_data1[887]), .S(n4265), .Z(
        n9180) );
  CMXI2X1 U18796 ( .A0(n9180), .A1(n9174), .S(n4017), .Z(n9187) );
  CMX2X1 U18797 ( .A0(n9175), .A1(n9187), .S(n4360), .Z(n9204) );
  CMXI2X1 U18798 ( .A0(n9176), .A1(n9204), .S(n3326), .Z(N2948) );
  CMX2X1 U18799 ( .A0(mem_data1[887]), .A1(mem_data1[888]), .S(n4265), .Z(
        n9183) );
  CMXI2X1 U18800 ( .A0(n9183), .A1(n9177), .S(n4017), .Z(n9190) );
  CMX2X1 U18801 ( .A0(n9178), .A1(n9190), .S(n3771), .Z(n9207) );
  CMXI2X1 U18802 ( .A0(n9179), .A1(n9207), .S(n3326), .Z(N2949) );
  CMX2X1 U18803 ( .A0(mem_data1[888]), .A1(mem_data1[889]), .S(n4265), .Z(
        n9186) );
  CMXI2X1 U18804 ( .A0(n9186), .A1(n9180), .S(n4017), .Z(n9193) );
  CMX2X1 U18805 ( .A0(n9181), .A1(n9193), .S(n3772), .Z(n9210) );
  CMXI2X1 U18806 ( .A0(n9182), .A1(n9210), .S(n3326), .Z(N2950) );
  CMX2X1 U18807 ( .A0(mem_data1[889]), .A1(mem_data1[890]), .S(n4265), .Z(
        n9189) );
  CMXI2X1 U18808 ( .A0(n9189), .A1(n9183), .S(n4017), .Z(n9196) );
  CMX2X1 U18809 ( .A0(n9184), .A1(n9196), .S(n3773), .Z(n9213) );
  CMXI2X1 U18810 ( .A0(n9185), .A1(n9213), .S(n3326), .Z(N2951) );
  CMX2X1 U18811 ( .A0(mem_data1[890]), .A1(mem_data1[891]), .S(n4265), .Z(
        n9192) );
  CMXI2X1 U18812 ( .A0(n9192), .A1(n9186), .S(n4017), .Z(n9203) );
  CMX2X1 U18813 ( .A0(n9187), .A1(n9203), .S(n3774), .Z(n9216) );
  CMXI2X1 U18814 ( .A0(n9188), .A1(n9216), .S(n3326), .Z(N2952) );
  CMX2X1 U18815 ( .A0(mem_data1[891]), .A1(mem_data1[892]), .S(n4265), .Z(
        n9195) );
  CMXI2X1 U18816 ( .A0(n9195), .A1(n9189), .S(n4017), .Z(n9206) );
  CMX2X1 U18817 ( .A0(n9190), .A1(n9206), .S(n3775), .Z(n9219) );
  CMXI2X1 U18818 ( .A0(n9191), .A1(n9219), .S(n3325), .Z(N2953) );
  CMX2X1 U18819 ( .A0(mem_data1[892]), .A1(mem_data1[893]), .S(n4265), .Z(
        n9202) );
  CMXI2X1 U18820 ( .A0(n9202), .A1(n9192), .S(n4017), .Z(n9209) );
  CMX2X1 U18821 ( .A0(n9193), .A1(n9209), .S(n3776), .Z(n9222) );
  CMXI2X1 U18822 ( .A0(n9194), .A1(n9222), .S(n3325), .Z(N2954) );
  CMX2X1 U18823 ( .A0(mem_data1[893]), .A1(mem_data1[894]), .S(n4265), .Z(
        n9205) );
  CMXI2X1 U18824 ( .A0(n9205), .A1(n9195), .S(n4017), .Z(n9212) );
  CMX2X1 U18825 ( .A0(n9196), .A1(n9212), .S(n3777), .Z(n9225) );
  CMXI2X1 U18826 ( .A0(n9197), .A1(n9225), .S(n3325), .Z(N2955) );
  CMXI2X1 U18827 ( .A0(n9199), .A1(n9198), .S(n4017), .Z(n9334) );
  CMX2X1 U18828 ( .A0(n9200), .A1(n9334), .S(n3790), .Z(n9463) );
  CMXI2X1 U18829 ( .A0(n9201), .A1(n9463), .S(n3328), .Z(N2163) );
  CMX2X1 U18830 ( .A0(mem_data1[894]), .A1(mem_data1[895]), .S(n4265), .Z(
        n9208) );
  CMXI2X1 U18831 ( .A0(n9208), .A1(n9202), .S(n4017), .Z(n9215) );
  CMX2X1 U18832 ( .A0(n9203), .A1(n9215), .S(n3791), .Z(n9228) );
  CMXI2X1 U18833 ( .A0(n9204), .A1(n9228), .S(n3328), .Z(N2956) );
  CMX2X1 U18834 ( .A0(mem_data1[895]), .A1(mem_data1[896]), .S(n4265), .Z(
        n9211) );
  CMXI2X1 U18835 ( .A0(n9211), .A1(n9205), .S(n4017), .Z(n9218) );
  CMX2X1 U18836 ( .A0(n9206), .A1(n9218), .S(n3812), .Z(n9231) );
  CMXI2X1 U18837 ( .A0(n9207), .A1(n9231), .S(n3328), .Z(N2957) );
  CMX2X1 U18838 ( .A0(mem_data1[896]), .A1(mem_data1[897]), .S(n4265), .Z(
        n9214) );
  CMXI2X1 U18839 ( .A0(n9214), .A1(n9208), .S(n4017), .Z(n9221) );
  CMX2X1 U18840 ( .A0(n9209), .A1(n9221), .S(n3811), .Z(n9237) );
  CMXI2X1 U18841 ( .A0(n9210), .A1(n9237), .S(n3328), .Z(N2958) );
  CMX2X1 U18842 ( .A0(mem_data1[897]), .A1(mem_data1[898]), .S(n4264), .Z(
        n9217) );
  CMXI2X1 U18843 ( .A0(n9217), .A1(n9211), .S(n4017), .Z(n9224) );
  CMX2X1 U18844 ( .A0(n9212), .A1(n9224), .S(n3790), .Z(n9240) );
  CMXI2X1 U18845 ( .A0(n9213), .A1(n9240), .S(n3328), .Z(N2959) );
  CMX2X1 U18846 ( .A0(mem_data1[898]), .A1(mem_data1[899]), .S(n4264), .Z(
        n9220) );
  CMXI2X1 U18847 ( .A0(n9220), .A1(n9214), .S(n4016), .Z(n9227) );
  CMX2X1 U18848 ( .A0(n9215), .A1(n9227), .S(n3791), .Z(n9243) );
  CMXI2X1 U18849 ( .A0(n9216), .A1(n9243), .S(n3328), .Z(N2960) );
  CMX2X1 U18850 ( .A0(mem_data1[899]), .A1(mem_data1[900]), .S(n4264), .Z(
        n9223) );
  CMXI2X1 U18851 ( .A0(n9223), .A1(n9217), .S(n4016), .Z(n9230) );
  CMX2X1 U18852 ( .A0(n9218), .A1(n9230), .S(n3792), .Z(n9246) );
  CMXI2X1 U18853 ( .A0(n9219), .A1(n9246), .S(n3328), .Z(N2961) );
  CMX2X1 U18854 ( .A0(mem_data1[900]), .A1(mem_data1[901]), .S(n4264), .Z(
        n9226) );
  CMXI2X1 U18855 ( .A0(n9226), .A1(n9220), .S(n4016), .Z(n9236) );
  CMX2X1 U18856 ( .A0(n9221), .A1(n9236), .S(n3793), .Z(n9249) );
  CMXI2X1 U18857 ( .A0(n9222), .A1(n9249), .S(n3328), .Z(N2962) );
  CMX2X1 U18858 ( .A0(mem_data1[901]), .A1(mem_data1[902]), .S(n4264), .Z(
        n9229) );
  CMXI2X1 U18859 ( .A0(n9229), .A1(n9223), .S(n4016), .Z(n9239) );
  CMX2X1 U18860 ( .A0(n9224), .A1(n9239), .S(n3794), .Z(n9252) );
  CMXI2X1 U18861 ( .A0(n9225), .A1(n9252), .S(n3328), .Z(N2963) );
  CMX2X1 U18862 ( .A0(mem_data1[902]), .A1(mem_data1[903]), .S(n4264), .Z(
        n9235) );
  CMXI2X1 U18863 ( .A0(n9235), .A1(n9226), .S(n4016), .Z(n9242) );
  CMX2X1 U18864 ( .A0(n9227), .A1(n9242), .S(n3792), .Z(n9255) );
  CMXI2X1 U18865 ( .A0(n9228), .A1(n9255), .S(n3328), .Z(N2964) );
  CMX2X1 U18866 ( .A0(mem_data1[903]), .A1(mem_data1[904]), .S(n4264), .Z(
        n9238) );
  CMXI2X1 U18867 ( .A0(n9238), .A1(n9229), .S(n4016), .Z(n9245) );
  CMX2X1 U18868 ( .A0(n9230), .A1(n9245), .S(n3792), .Z(n9258) );
  CMXI2X1 U18869 ( .A0(n9231), .A1(n9258), .S(n3328), .Z(N2965) );
  CMX2X1 U18870 ( .A0(n9233), .A1(n9232), .S(n3793), .Z(n9495) );
  CMXI2X1 U18871 ( .A0(n9234), .A1(n9495), .S(n3327), .Z(N2164) );
  CMX2X1 U18872 ( .A0(mem_data1[904]), .A1(mem_data1[905]), .S(n4264), .Z(
        n9241) );
  CMXI2X1 U18873 ( .A0(n9241), .A1(n9235), .S(n4016), .Z(n9248) );
  CMX2X1 U18874 ( .A0(n9236), .A1(n9248), .S(n3794), .Z(n9261) );
  CMXI2X1 U18875 ( .A0(n9237), .A1(n9261), .S(n3327), .Z(N2966) );
  CMX2X1 U18876 ( .A0(mem_data1[905]), .A1(mem_data1[906]), .S(n4264), .Z(
        n9244) );
  CMXI2X1 U18877 ( .A0(n9244), .A1(n9238), .S(n4016), .Z(n9251) );
  CMX2X1 U18878 ( .A0(n9239), .A1(n9251), .S(n3795), .Z(n9264) );
  CMXI2X1 U18879 ( .A0(n9240), .A1(n9264), .S(n3327), .Z(N2967) );
  CMX2X1 U18880 ( .A0(mem_data1[906]), .A1(mem_data1[907]), .S(n4264), .Z(
        n9247) );
  CMXI2X1 U18881 ( .A0(n9247), .A1(n9241), .S(n4016), .Z(n9254) );
  CMX2X1 U18882 ( .A0(n9242), .A1(n9254), .S(n3796), .Z(n9272) );
  CMXI2X1 U18883 ( .A0(n9243), .A1(n9272), .S(n3327), .Z(N2968) );
  CMX2X1 U18884 ( .A0(mem_data1[907]), .A1(mem_data1[908]), .S(n4264), .Z(
        n9250) );
  CMXI2X1 U18885 ( .A0(n9250), .A1(n9244), .S(n4016), .Z(n9257) );
  CMX2X1 U18886 ( .A0(n9245), .A1(n9257), .S(n3797), .Z(n9275) );
  CMXI2X1 U18887 ( .A0(n9246), .A1(n9275), .S(n3327), .Z(N2969) );
  CMX2X1 U18888 ( .A0(mem_data1[908]), .A1(mem_data1[909]), .S(n4263), .Z(
        n9253) );
  CMXI2X1 U18889 ( .A0(n9253), .A1(n9247), .S(n4016), .Z(n9260) );
  CMX2X1 U18890 ( .A0(n9248), .A1(n9260), .S(n3805), .Z(n9278) );
  CMXI2X1 U18891 ( .A0(n9249), .A1(n9278), .S(n3327), .Z(N2970) );
  CMX2X1 U18892 ( .A0(mem_data1[909]), .A1(mem_data1[910]), .S(n4263), .Z(
        n9256) );
  CMXI2X1 U18893 ( .A0(n9256), .A1(n9250), .S(n4016), .Z(n9263) );
  CMX2X1 U18894 ( .A0(n9251), .A1(n9263), .S(n3806), .Z(n9281) );
  CMXI2X1 U18895 ( .A0(n9252), .A1(n9281), .S(n3327), .Z(N2971) );
  CMX2X1 U18896 ( .A0(mem_data1[910]), .A1(mem_data1[911]), .S(n4263), .Z(
        n9259) );
  CMXI2X1 U18897 ( .A0(n9259), .A1(n9253), .S(n4016), .Z(n9271) );
  CMX2X1 U18898 ( .A0(n9254), .A1(n9271), .S(n3807), .Z(n9284) );
  CMXI2X1 U18899 ( .A0(n9255), .A1(n9284), .S(n3330), .Z(N2972) );
  CMX2X1 U18900 ( .A0(mem_data1[911]), .A1(mem_data1[912]), .S(n4263), .Z(
        n9262) );
  CMXI2X1 U18901 ( .A0(n9262), .A1(n9256), .S(n4016), .Z(n9274) );
  CMX2X1 U18902 ( .A0(n9257), .A1(n9274), .S(n3808), .Z(n9287) );
  CMXI2X1 U18903 ( .A0(n9258), .A1(n9287), .S(n3330), .Z(N2973) );
  CMX2X1 U18904 ( .A0(mem_data1[912]), .A1(mem_data1[913]), .S(n4263), .Z(
        n9270) );
  CMXI2X1 U18905 ( .A0(n9270), .A1(n9259), .S(n4016), .Z(n9277) );
  CMX2X1 U18906 ( .A0(n9260), .A1(n9277), .S(n3809), .Z(n9290) );
  CMXI2X1 U18907 ( .A0(n9261), .A1(n9290), .S(n3330), .Z(N2974) );
  CMX2X1 U18908 ( .A0(mem_data1[913]), .A1(mem_data1[914]), .S(n4263), .Z(
        n9273) );
  CMXI2X1 U18909 ( .A0(n9273), .A1(n9262), .S(n4016), .Z(n9280) );
  CMX2X1 U18910 ( .A0(n9263), .A1(n9280), .S(n3810), .Z(n9293) );
  CMXI2X1 U18911 ( .A0(n9264), .A1(n9293), .S(n3330), .Z(N2975) );
  CMX2X1 U18912 ( .A0(n9266), .A1(n9265), .S(n3811), .Z(n9527) );
  CMXI2X1 U18913 ( .A0(n9267), .A1(n9527), .S(n3330), .Z(N2165) );
  CMXI2X1 U18914 ( .A0(n9269), .A1(n9268), .S(n3330), .Z(N2084) );
  CMX2X1 U18915 ( .A0(mem_data1[914]), .A1(mem_data1[915]), .S(n4263), .Z(
        n9276) );
  CMXI2X1 U18916 ( .A0(n9276), .A1(n9270), .S(n4015), .Z(n9283) );
  CMX2X1 U18917 ( .A0(n9271), .A1(n9283), .S(n3812), .Z(n9296) );
  CMXI2X1 U18918 ( .A0(n9272), .A1(n9296), .S(n3330), .Z(N2976) );
  CMX2X1 U18919 ( .A0(mem_data1[915]), .A1(mem_data1[916]), .S(n4263), .Z(
        n9279) );
  CMXI2X1 U18920 ( .A0(n9279), .A1(n9273), .S(n4015), .Z(n9286) );
  CMX2X1 U18921 ( .A0(n9274), .A1(n9286), .S(n4363), .Z(n9299) );
  CMXI2X1 U18922 ( .A0(n9275), .A1(n9299), .S(n3329), .Z(N2977) );
  CMX2X1 U18923 ( .A0(mem_data1[916]), .A1(mem_data1[917]), .S(n4263), .Z(
        n9282) );
  CMXI2X1 U18924 ( .A0(n9282), .A1(n9276), .S(n4015), .Z(n9289) );
  CMX2X1 U18925 ( .A0(n9277), .A1(n9289), .S(n3771), .Z(n9305) );
  CMXI2X1 U18926 ( .A0(n9278), .A1(n9305), .S(n3329), .Z(N2978) );
  CMX2X1 U18927 ( .A0(mem_data1[917]), .A1(mem_data1[918]), .S(n4263), .Z(
        n9285) );
  CMXI2X1 U18928 ( .A0(n9285), .A1(n9279), .S(n4015), .Z(n9292) );
  CMX2X1 U18929 ( .A0(n9280), .A1(n9292), .S(n4367), .Z(n9308) );
  CMXI2X1 U18930 ( .A0(n9281), .A1(n9308), .S(n3329), .Z(N2979) );
  CMX2X1 U18931 ( .A0(mem_data1[918]), .A1(mem_data1[919]), .S(n4263), .Z(
        n9288) );
  CMXI2X1 U18932 ( .A0(n9288), .A1(n9282), .S(n4015), .Z(n9295) );
  CMX2X1 U18933 ( .A0(n9283), .A1(n9295), .S(n3812), .Z(n9311) );
  CMXI2X1 U18934 ( .A0(n9284), .A1(n9311), .S(n3329), .Z(N2980) );
  CMX2X1 U18935 ( .A0(mem_data1[919]), .A1(mem_data1[920]), .S(n4262), .Z(
        n9291) );
  CMXI2X1 U18936 ( .A0(n9291), .A1(n9285), .S(n4015), .Z(n9298) );
  CMX2X1 U18937 ( .A0(n9286), .A1(n9298), .S(n3795), .Z(n9314) );
  CMXI2X1 U18938 ( .A0(n9287), .A1(n9314), .S(n3329), .Z(N2981) );
  CMX2X1 U18939 ( .A0(mem_data1[920]), .A1(mem_data1[921]), .S(n4262), .Z(
        n9294) );
  CMXI2X1 U18940 ( .A0(n9294), .A1(n9288), .S(n4015), .Z(n9304) );
  CMX2X1 U18941 ( .A0(n9289), .A1(n9304), .S(n3796), .Z(n9317) );
  CMXI2X1 U18942 ( .A0(n9290), .A1(n9317), .S(n3329), .Z(N2982) );
  CMX2X1 U18943 ( .A0(mem_data1[921]), .A1(mem_data1[922]), .S(n4262), .Z(
        n9297) );
  CMXI2X1 U18944 ( .A0(n9297), .A1(n9291), .S(n4015), .Z(n9307) );
  CMX2X1 U18945 ( .A0(n9292), .A1(n9307), .S(n3797), .Z(n9320) );
  CMXI2X1 U18946 ( .A0(n9293), .A1(n9320), .S(n3329), .Z(N2983) );
  CMX2X1 U18947 ( .A0(mem_data1[922]), .A1(mem_data1[923]), .S(n4262), .Z(
        n9303) );
  CMXI2X1 U18948 ( .A0(n9303), .A1(n9294), .S(n4015), .Z(n9310) );
  CMX2X1 U18949 ( .A0(n9295), .A1(n9310), .S(n3805), .Z(n9323) );
  CMXI2X1 U18950 ( .A0(n9296), .A1(n9323), .S(n3329), .Z(N2984) );
  CMX2X1 U18951 ( .A0(mem_data1[923]), .A1(mem_data1[924]), .S(n4262), .Z(
        n9306) );
  CMXI2X1 U18952 ( .A0(n9306), .A1(n9297), .S(n4015), .Z(n9313) );
  CMX2X1 U18953 ( .A0(n9298), .A1(n9313), .S(n3806), .Z(n9326) );
  CMXI2X1 U18954 ( .A0(n9299), .A1(n9326), .S(n3329), .Z(N2985) );
  CMX2X1 U18955 ( .A0(n9301), .A1(n9300), .S(n3793), .Z(n9561) );
  CMXI2X1 U18956 ( .A0(n9302), .A1(n9561), .S(n3329), .Z(N2166) );
  CMX2X1 U18957 ( .A0(mem_data1[924]), .A1(mem_data1[925]), .S(n4262), .Z(
        n9309) );
  CMXI2X1 U18958 ( .A0(n9309), .A1(n9303), .S(n4015), .Z(n9316) );
  CMX2X1 U18959 ( .A0(n9304), .A1(n9316), .S(n3772), .Z(n9329) );
  CMXI2X1 U18960 ( .A0(n9305), .A1(n9329), .S(n3329), .Z(N2986) );
  CMX2X1 U18961 ( .A0(mem_data1[925]), .A1(mem_data1[926]), .S(n4262), .Z(
        n9312) );
  CMXI2X1 U18962 ( .A0(n9312), .A1(n9306), .S(n4015), .Z(n9319) );
  CMX2X1 U18963 ( .A0(n9307), .A1(n9319), .S(n3773), .Z(n9332) );
  CMXI2X1 U18964 ( .A0(n9308), .A1(n9332), .S(n3332), .Z(N2987) );
  CMX2X1 U18965 ( .A0(mem_data1[926]), .A1(mem_data1[927]), .S(n4262), .Z(
        n9315) );
  CMXI2X1 U18966 ( .A0(n9315), .A1(n9309), .S(n4015), .Z(n9322) );
  CMX2X1 U18967 ( .A0(n9310), .A1(n9322), .S(n3774), .Z(n9338) );
  CMXI2X1 U18968 ( .A0(n9311), .A1(n9338), .S(n3332), .Z(N2988) );
  CMX2X1 U18969 ( .A0(mem_data1[927]), .A1(mem_data1[928]), .S(n4262), .Z(
        n9318) );
  CMXI2X1 U18970 ( .A0(n9318), .A1(n9312), .S(n4015), .Z(n9325) );
  CMX2X1 U18971 ( .A0(n9313), .A1(n9325), .S(n3775), .Z(n9341) );
  CMXI2X1 U18972 ( .A0(n9314), .A1(n9341), .S(n3332), .Z(N2989) );
  CMX2X1 U18973 ( .A0(mem_data1[928]), .A1(mem_data1[929]), .S(n4262), .Z(
        n9321) );
  CMXI2X1 U18974 ( .A0(n9321), .A1(n9315), .S(n4015), .Z(n9328) );
  CMX2X1 U18975 ( .A0(n9316), .A1(n9328), .S(n3776), .Z(n9344) );
  CMXI2X1 U18976 ( .A0(n9317), .A1(n9344), .S(n3331), .Z(N2990) );
  CMX2X1 U18977 ( .A0(mem_data1[929]), .A1(mem_data1[930]), .S(n4262), .Z(
        n9324) );
  CMXI2X1 U18978 ( .A0(n9324), .A1(n9318), .S(n4015), .Z(n9331) );
  CMX2X1 U18979 ( .A0(n9319), .A1(n9331), .S(n3777), .Z(n9347) );
  CMXI2X1 U18980 ( .A0(n9320), .A1(n9347), .S(n3331), .Z(N2991) );
  CMX2X1 U18981 ( .A0(mem_data1[930]), .A1(mem_data1[931]), .S(n4261), .Z(
        n9327) );
  CMXI2X1 U18982 ( .A0(n9327), .A1(n9321), .S(n4014), .Z(n9337) );
  CMX2X1 U18983 ( .A0(n9322), .A1(n9337), .S(n3790), .Z(n9350) );
  CMXI2X1 U18984 ( .A0(n9323), .A1(n9350), .S(n3331), .Z(N2992) );
  CMX2X1 U18985 ( .A0(mem_data1[931]), .A1(mem_data1[932]), .S(n4261), .Z(
        n9330) );
  CMXI2X1 U18986 ( .A0(n9330), .A1(n9324), .S(n4014), .Z(n9340) );
  CMX2X1 U18987 ( .A0(n9325), .A1(n9340), .S(n3791), .Z(n9353) );
  CMXI2X1 U18988 ( .A0(n9326), .A1(n9353), .S(n3331), .Z(N2993) );
  CMX2X1 U18989 ( .A0(mem_data1[932]), .A1(mem_data1[933]), .S(n4261), .Z(
        n9336) );
  CMXI2X1 U18990 ( .A0(n9336), .A1(n9327), .S(n4014), .Z(n9343) );
  CMX2X1 U18991 ( .A0(n9328), .A1(n9343), .S(n3792), .Z(n9356) );
  CMXI2X1 U18992 ( .A0(n9329), .A1(n9356), .S(n3331), .Z(N2994) );
  CMX2X1 U18993 ( .A0(mem_data1[933]), .A1(mem_data1[934]), .S(n4261), .Z(
        n9339) );
  CMXI2X1 U18994 ( .A0(n9339), .A1(n9330), .S(n4014), .Z(n9346) );
  CMX2X1 U18995 ( .A0(n9331), .A1(n9346), .S(n3793), .Z(n9359) );
  CMXI2X1 U18996 ( .A0(n9332), .A1(n9359), .S(n3331), .Z(N2995) );
  CMX2X1 U18997 ( .A0(n9334), .A1(n9333), .S(n3794), .Z(n9585) );
  CMXI2X1 U18998 ( .A0(n9335), .A1(n9585), .S(n3331), .Z(N2167) );
  CMX2X1 U18999 ( .A0(mem_data1[934]), .A1(mem_data1[935]), .S(n4261), .Z(
        n9342) );
  CMXI2X1 U19000 ( .A0(n9342), .A1(n9336), .S(n4014), .Z(n9349) );
  CMX2X1 U19001 ( .A0(n9337), .A1(n9349), .S(n3795), .Z(n9362) );
  CMXI2X1 U19002 ( .A0(n9338), .A1(n9362), .S(n3331), .Z(N2996) );
  CMX2X1 U19003 ( .A0(mem_data1[935]), .A1(mem_data1[936]), .S(n4261), .Z(
        n9345) );
  CMXI2X1 U19004 ( .A0(n9345), .A1(n9339), .S(n4014), .Z(n9352) );
  CMX2X1 U19005 ( .A0(n9340), .A1(n9352), .S(n3796), .Z(n9365) );
  CMXI2X1 U19006 ( .A0(n9341), .A1(n9365), .S(n3331), .Z(N2997) );
  CMX2X1 U19007 ( .A0(mem_data1[936]), .A1(mem_data1[937]), .S(n4270), .Z(
        n9348) );
  CMXI2X1 U19008 ( .A0(n9348), .A1(n9342), .S(n4014), .Z(n9355) );
  CMX2X1 U19009 ( .A0(n9343), .A1(n9355), .S(n3797), .Z(n9370) );
  CMXI2X1 U19010 ( .A0(n9344), .A1(n9370), .S(n3331), .Z(N2998) );
  CMX2X1 U19011 ( .A0(mem_data1[937]), .A1(mem_data1[938]), .S(n4293), .Z(
        n9351) );
  CMXI2X1 U19012 ( .A0(n9351), .A1(n9345), .S(n4014), .Z(n9358) );
  CMX2X1 U19013 ( .A0(n9346), .A1(n9358), .S(n3805), .Z(n9373) );
  CMXI2X1 U19014 ( .A0(n9347), .A1(n9373), .S(n3331), .Z(N2999) );
  CMX2X1 U19015 ( .A0(mem_data1[938]), .A1(mem_data1[939]), .S(n4293), .Z(
        n9354) );
  CMXI2X1 U19016 ( .A0(n9354), .A1(n9348), .S(n4014), .Z(n9361) );
  CMX2X1 U19017 ( .A0(n9349), .A1(n9361), .S(n3806), .Z(n9376) );
  CMXI2X1 U19018 ( .A0(n9350), .A1(n9376), .S(n3330), .Z(N3000) );
  CMX2X1 U19019 ( .A0(mem_data1[939]), .A1(mem_data1[940]), .S(n4293), .Z(
        n9357) );
  CMXI2X1 U19020 ( .A0(n9357), .A1(n9351), .S(n4014), .Z(n9364) );
  CMX2X1 U19021 ( .A0(n9352), .A1(n9364), .S(n3771), .Z(n9379) );
  CMXI2X1 U19022 ( .A0(n9353), .A1(n9379), .S(n3330), .Z(N3001) );
  CMX2X1 U19023 ( .A0(mem_data1[940]), .A1(mem_data1[941]), .S(n4293), .Z(
        n9360) );
  CMXI2X1 U19024 ( .A0(n9360), .A1(n9354), .S(n4014), .Z(n9369) );
  CMX2X1 U19025 ( .A0(n9355), .A1(n9369), .S(n4359), .Z(n9382) );
  CMXI2X1 U19026 ( .A0(n9356), .A1(n9382), .S(n3330), .Z(N3002) );
  CMX2X1 U19027 ( .A0(mem_data1[941]), .A1(mem_data1[942]), .S(n4293), .Z(
        n9363) );
  CMXI2X1 U19028 ( .A0(n9363), .A1(n9357), .S(n4014), .Z(n9372) );
  CMX2X1 U19029 ( .A0(n9358), .A1(n9372), .S(n3807), .Z(n9385) );
  CMXI2X1 U19030 ( .A0(n9359), .A1(n9385), .S(n3330), .Z(N3003) );
  CMX2X1 U19031 ( .A0(mem_data1[942]), .A1(mem_data1[943]), .S(n4293), .Z(
        n9368) );
  CMXI2X1 U19032 ( .A0(n9368), .A1(n9360), .S(n4014), .Z(n9375) );
  CMX2X1 U19033 ( .A0(n9361), .A1(n9375), .S(n3796), .Z(n9388) );
  CMXI2X1 U19034 ( .A0(n9362), .A1(n9388), .S(n3299), .Z(N3004) );
  CMX2X1 U19035 ( .A0(mem_data1[943]), .A1(mem_data1[944]), .S(n4293), .Z(
        n9371) );
  CMXI2X1 U19036 ( .A0(n9371), .A1(n9363), .S(n4014), .Z(n9378) );
  CMX2X1 U19037 ( .A0(n9364), .A1(n9378), .S(n3805), .Z(n9391) );
  CMXI2X1 U19038 ( .A0(n9365), .A1(n9391), .S(n3299), .Z(N3005) );
  CMXI2X1 U19039 ( .A0(n9367), .A1(n9366), .S(n3299), .Z(N2168) );
  CMX2X1 U19040 ( .A0(mem_data1[944]), .A1(mem_data1[945]), .S(n4293), .Z(
        n9374) );
  CMXI2X1 U19041 ( .A0(n9374), .A1(n9368), .S(n4014), .Z(n9381) );
  CMX2X1 U19042 ( .A0(n9369), .A1(n9381), .S(n3806), .Z(n9394) );
  CMXI2X1 U19043 ( .A0(n9370), .A1(n9394), .S(n3299), .Z(N3006) );
  CMX2X1 U19044 ( .A0(mem_data1[945]), .A1(mem_data1[946]), .S(n4293), .Z(
        n9377) );
  CMXI2X1 U19045 ( .A0(n9377), .A1(n9371), .S(n4014), .Z(n9384) );
  CMX2X1 U19046 ( .A0(n9372), .A1(n9384), .S(n3777), .Z(n9397) );
  CMXI2X1 U19047 ( .A0(n9373), .A1(n9397), .S(n3299), .Z(N3007) );
  CMX2X1 U19048 ( .A0(mem_data1[946]), .A1(mem_data1[947]), .S(n4293), .Z(
        n9380) );
  CMXI2X1 U19049 ( .A0(n9380), .A1(n9374), .S(n4013), .Z(n9387) );
  CMX2X1 U19050 ( .A0(n9375), .A1(n9387), .S(n3790), .Z(n9402) );
  CMXI2X1 U19051 ( .A0(n9376), .A1(n9402), .S(n3477), .Z(N3008) );
  CMX2X1 U19052 ( .A0(mem_data1[947]), .A1(mem_data1[948]), .S(n4238), .Z(
        n9383) );
  CMXI2X1 U19053 ( .A0(n9383), .A1(n9377), .S(n4013), .Z(n9390) );
  CMX2X1 U19054 ( .A0(n9378), .A1(n9390), .S(n3791), .Z(n9405) );
  CMXI2X1 U19055 ( .A0(n9379), .A1(n9405), .S(n3476), .Z(N3009) );
  CMX2X1 U19056 ( .A0(mem_data1[948]), .A1(mem_data1[949]), .S(n4238), .Z(
        n9386) );
  CMXI2X1 U19057 ( .A0(n9386), .A1(n9380), .S(n4013), .Z(n9393) );
  CMX2X1 U19058 ( .A0(n9381), .A1(n9393), .S(n3792), .Z(n9408) );
  CMXI2X1 U19059 ( .A0(n9382), .A1(n9408), .S(n3475), .Z(N3010) );
  CMX2X1 U19060 ( .A0(mem_data1[949]), .A1(mem_data1[950]), .S(n4237), .Z(
        n9389) );
  CMXI2X1 U19061 ( .A0(n9389), .A1(n9383), .S(n4013), .Z(n9396) );
  CMX2X1 U19062 ( .A0(n9384), .A1(n9396), .S(n3793), .Z(n9411) );
  CMXI2X1 U19063 ( .A0(n9385), .A1(n9411), .S(n3474), .Z(N3011) );
  CMX2X1 U19064 ( .A0(mem_data1[950]), .A1(mem_data1[951]), .S(n4238), .Z(
        n9392) );
  CMXI2X1 U19065 ( .A0(n9392), .A1(n9386), .S(n4013), .Z(n9401) );
  CMX2X1 U19066 ( .A0(n9387), .A1(n9401), .S(n3775), .Z(n9414) );
  CMXI2X1 U19067 ( .A0(n9388), .A1(n9414), .S(n3473), .Z(N3012) );
  CMX2X1 U19068 ( .A0(mem_data1[951]), .A1(mem_data1[952]), .S(n4237), .Z(
        n9395) );
  CMXI2X1 U19069 ( .A0(n9395), .A1(n9389), .S(n4013), .Z(n9404) );
  CMX2X1 U19070 ( .A0(n9390), .A1(n9404), .S(n3772), .Z(n9417) );
  CMXI2X1 U19071 ( .A0(n9391), .A1(n9417), .S(n3472), .Z(N3013) );
  CMX2X1 U19072 ( .A0(mem_data1[952]), .A1(mem_data1[953]), .S(n4238), .Z(
        n9400) );
  CMXI2X1 U19073 ( .A0(n9400), .A1(n9392), .S(n4013), .Z(n9407) );
  CMX2X1 U19074 ( .A0(n9393), .A1(n9407), .S(n3773), .Z(n9420) );
  CMXI2X1 U19075 ( .A0(n9394), .A1(n9420), .S(n3285), .Z(N3014) );
  CMX2X1 U19076 ( .A0(mem_data1[953]), .A1(mem_data1[954]), .S(n4237), .Z(
        n9403) );
  CMXI2X1 U19077 ( .A0(n9403), .A1(n9395), .S(n4013), .Z(n9410) );
  CMX2X1 U19078 ( .A0(n9396), .A1(n9410), .S(n3774), .Z(n9423) );
  CMXI2X1 U19079 ( .A0(n9397), .A1(n9423), .S(n3285), .Z(N3015) );
  CMXI2X1 U19080 ( .A0(n9399), .A1(n9398), .S(n3285), .Z(N2169) );
  CMX2X1 U19081 ( .A0(mem_data1[954]), .A1(mem_data1[955]), .S(n4238), .Z(
        n9406) );
  CMXI2X1 U19082 ( .A0(n9406), .A1(n9400), .S(n4013), .Z(n9413) );
  CMX2X1 U19083 ( .A0(n9401), .A1(n9413), .S(n3775), .Z(n9426) );
  CMXI2X1 U19084 ( .A0(n9402), .A1(n9426), .S(n3285), .Z(N3016) );
  CMX2X1 U19085 ( .A0(mem_data1[955]), .A1(mem_data1[956]), .S(n4237), .Z(
        n9409) );
  CMXI2X1 U19086 ( .A0(n9409), .A1(n9403), .S(n4013), .Z(n9416) );
  CMX2X1 U19087 ( .A0(n9404), .A1(n9416), .S(n3805), .Z(n9429) );
  CMXI2X1 U19088 ( .A0(n9405), .A1(n9429), .S(n3285), .Z(N3017) );
  CMX2X1 U19089 ( .A0(mem_data1[956]), .A1(mem_data1[957]), .S(n4238), .Z(
        n9412) );
  CMXI2X1 U19090 ( .A0(n9412), .A1(n9406), .S(n4013), .Z(n9419) );
  CMX2X1 U19091 ( .A0(n9407), .A1(n9419), .S(n3806), .Z(n9434) );
  CMXI2X1 U19092 ( .A0(n9408), .A1(n9434), .S(n3285), .Z(N3018) );
  CMX2X1 U19093 ( .A0(mem_data1[957]), .A1(mem_data1[958]), .S(n4237), .Z(
        n9415) );
  CMXI2X1 U19094 ( .A0(n9415), .A1(n9409), .S(n4013), .Z(n9422) );
  CMX2X1 U19095 ( .A0(n9410), .A1(n9422), .S(n3777), .Z(n9437) );
  CMXI2X1 U19096 ( .A0(n9411), .A1(n9437), .S(n3441), .Z(N3019) );
  CMX2X1 U19097 ( .A0(mem_data1[958]), .A1(mem_data1[959]), .S(n4292), .Z(
        n9418) );
  CMXI2X1 U19098 ( .A0(n9418), .A1(n9412), .S(n4013), .Z(n9425) );
  CMX2X1 U19099 ( .A0(n9413), .A1(n9425), .S(n3776), .Z(n9440) );
  CMXI2X1 U19100 ( .A0(n9414), .A1(n9440), .S(n3443), .Z(N3020) );
  CMX2X1 U19101 ( .A0(mem_data1[959]), .A1(mem_data1[960]), .S(n4292), .Z(
        n9421) );
  CMXI2X1 U19102 ( .A0(n9421), .A1(n9415), .S(n4013), .Z(n9428) );
  CMX2X1 U19103 ( .A0(n9416), .A1(n9428), .S(n4367), .Z(n9443) );
  CMXI2X1 U19104 ( .A0(n9417), .A1(n9443), .S(n3444), .Z(N3021) );
  CMX2X1 U19105 ( .A0(mem_data1[960]), .A1(mem_data1[961]), .S(n4292), .Z(
        n9424) );
  CMXI2X1 U19106 ( .A0(n9424), .A1(n9418), .S(n4013), .Z(n9433) );
  CMX2X1 U19107 ( .A0(n9419), .A1(n9433), .S(n3771), .Z(n9446) );
  CMXI2X1 U19108 ( .A0(n9420), .A1(n9446), .S(n3445), .Z(N3022) );
  CMX2X1 U19109 ( .A0(mem_data1[961]), .A1(mem_data1[962]), .S(n4292), .Z(
        n9427) );
  CMXI2X1 U19110 ( .A0(n9427), .A1(n9421), .S(n4013), .Z(n9436) );
  CMX2X1 U19111 ( .A0(n9422), .A1(n9436), .S(n3772), .Z(n9449) );
  CMXI2X1 U19112 ( .A0(n9423), .A1(n9449), .S(n3447), .Z(N3023) );
  CMX2X1 U19113 ( .A0(mem_data1[962]), .A1(mem_data1[963]), .S(n4292), .Z(
        n9432) );
  CMXI2X1 U19114 ( .A0(n9432), .A1(n9424), .S(n4012), .Z(n9439) );
  CMX2X1 U19115 ( .A0(n9425), .A1(n9439), .S(n3773), .Z(n9452) );
  CMXI2X1 U19116 ( .A0(n9426), .A1(n9452), .S(n3448), .Z(N3024) );
  CMX2X1 U19117 ( .A0(mem_data1[963]), .A1(mem_data1[964]), .S(n4292), .Z(
        n9435) );
  CMXI2X1 U19118 ( .A0(n9435), .A1(n9427), .S(n4012), .Z(n9442) );
  CMX2X1 U19119 ( .A0(n9428), .A1(n9442), .S(n3774), .Z(n9455) );
  CMXI2X1 U19120 ( .A0(n9429), .A1(n9455), .S(n3449), .Z(N3025) );
  CMXI2X1 U19121 ( .A0(n9431), .A1(n9430), .S(n3324), .Z(N2170) );
  CMX2X1 U19122 ( .A0(mem_data1[964]), .A1(mem_data1[965]), .S(n4292), .Z(
        n9438) );
  CMXI2X1 U19123 ( .A0(n9438), .A1(n9432), .S(n4012), .Z(n9445) );
  CMX2X1 U19124 ( .A0(n9433), .A1(n9445), .S(n3807), .Z(n9458) );
  CMXI2X1 U19125 ( .A0(n9434), .A1(n9458), .S(n3315), .Z(N3026) );
  CMX2X1 U19126 ( .A0(mem_data1[965]), .A1(mem_data1[966]), .S(n4292), .Z(
        n9441) );
  CMXI2X1 U19127 ( .A0(n9441), .A1(n9435), .S(n4012), .Z(n9448) );
  CMX2X1 U19128 ( .A0(n9436), .A1(n9448), .S(n3807), .Z(n9461) );
  CMXI2X1 U19129 ( .A0(n9437), .A1(n9461), .S(n3315), .Z(N3027) );
  CMX2X1 U19130 ( .A0(mem_data1[966]), .A1(mem_data1[967]), .S(n4292), .Z(
        n9444) );
  CMXI2X1 U19131 ( .A0(n9444), .A1(n9438), .S(n4012), .Z(n9451) );
  CMX2X1 U19132 ( .A0(n9439), .A1(n9451), .S(n3807), .Z(n9466) );
  CMXI2X1 U19133 ( .A0(n9440), .A1(n9466), .S(n3315), .Z(N3028) );
  CMX2X1 U19134 ( .A0(mem_data1[967]), .A1(mem_data1[968]), .S(n4292), .Z(
        n9447) );
  CMXI2X1 U19135 ( .A0(n9447), .A1(n9441), .S(n4012), .Z(n9454) );
  CMX2X1 U19136 ( .A0(n9442), .A1(n9454), .S(n3805), .Z(n9469) );
  CMXI2X1 U19137 ( .A0(n9443), .A1(n9469), .S(n3283), .Z(N3029) );
  CMX2X1 U19138 ( .A0(mem_data1[968]), .A1(mem_data1[969]), .S(n4292), .Z(
        n9450) );
  CMXI2X1 U19139 ( .A0(n9450), .A1(n9444), .S(n4012), .Z(n9457) );
  CMX2X1 U19140 ( .A0(n9445), .A1(n9457), .S(n3792), .Z(n9472) );
  CMXI2X1 U19141 ( .A0(n9446), .A1(n9472), .S(n3283), .Z(N3030) );
  CMX2X1 U19142 ( .A0(mem_data1[969]), .A1(mem_data1[970]), .S(n4291), .Z(
        n9453) );
  CMXI2X1 U19143 ( .A0(n9453), .A1(n9447), .S(n4012), .Z(n9460) );
  CMX2X1 U19144 ( .A0(n9448), .A1(n9460), .S(n3793), .Z(n9475) );
  CMXI2X1 U19145 ( .A0(n9449), .A1(n9475), .S(n3283), .Z(N3031) );
  CMX2X1 U19146 ( .A0(mem_data1[970]), .A1(mem_data1[971]), .S(n4291), .Z(
        n9456) );
  CMXI2X1 U19147 ( .A0(n9456), .A1(n9450), .S(n4012), .Z(n9465) );
  CMX2X1 U19148 ( .A0(n9451), .A1(n9465), .S(n3794), .Z(n9478) );
  CMXI2X1 U19149 ( .A0(n9452), .A1(n9478), .S(n3284), .Z(N3032) );
  CMX2X1 U19150 ( .A0(mem_data1[971]), .A1(mem_data1[972]), .S(n4291), .Z(
        n9459) );
  CMXI2X1 U19151 ( .A0(n9459), .A1(n9453), .S(n4012), .Z(n9468) );
  CMX2X1 U19152 ( .A0(n9454), .A1(n9468), .S(n3795), .Z(n9481) );
  CMXI2X1 U19153 ( .A0(n9455), .A1(n9481), .S(n3284), .Z(N3033) );
  CMX2X1 U19154 ( .A0(mem_data1[972]), .A1(mem_data1[973]), .S(n4291), .Z(
        n9464) );
  CMXI2X1 U19155 ( .A0(n9464), .A1(n9456), .S(n4012), .Z(n9471) );
  CMX2X1 U19156 ( .A0(n9457), .A1(n9471), .S(n3796), .Z(n9484) );
  CMXI2X1 U19157 ( .A0(n9458), .A1(n9484), .S(n3284), .Z(N3034) );
  CMX2X1 U19158 ( .A0(mem_data1[973]), .A1(mem_data1[974]), .S(n4291), .Z(
        n9467) );
  CMXI2X1 U19159 ( .A0(n9467), .A1(n9459), .S(n4012), .Z(n9474) );
  CMX2X1 U19160 ( .A0(n9460), .A1(n9474), .S(n3797), .Z(n9487) );
  CMXI2X1 U19161 ( .A0(n9461), .A1(n9487), .S(n3284), .Z(N3035) );
  CMXI2X1 U19162 ( .A0(n9463), .A1(n9462), .S(n3284), .Z(N2171) );
  CMX2X1 U19163 ( .A0(mem_data1[974]), .A1(mem_data1[975]), .S(n4291), .Z(
        n9470) );
  CMXI2X1 U19164 ( .A0(n9470), .A1(n9464), .S(n4012), .Z(n9477) );
  CMX2X1 U19165 ( .A0(n9465), .A1(n9477), .S(n3805), .Z(n9490) );
  CMXI2X1 U19166 ( .A0(n9466), .A1(n9490), .S(n3284), .Z(N3036) );
  CMX2X1 U19167 ( .A0(mem_data1[975]), .A1(mem_data1[976]), .S(n4291), .Z(
        n9473) );
  CMXI2X1 U19168 ( .A0(n9473), .A1(n9467), .S(n4012), .Z(n9480) );
  CMX2X1 U19169 ( .A0(n9468), .A1(n9480), .S(n3806), .Z(n9493) );
  CMXI2X1 U19170 ( .A0(n9469), .A1(n9493), .S(n3284), .Z(N3037) );
  CMX2X1 U19171 ( .A0(mem_data1[976]), .A1(mem_data1[977]), .S(n4291), .Z(
        n9476) );
  CMXI2X1 U19172 ( .A0(n9476), .A1(n9470), .S(n4012), .Z(n9483) );
  CMX2X1 U19173 ( .A0(n9471), .A1(n9483), .S(n3807), .Z(n9498) );
  CMXI2X1 U19174 ( .A0(n9472), .A1(n9498), .S(n3284), .Z(N3038) );
  CMX2X1 U19175 ( .A0(mem_data1[977]), .A1(mem_data1[978]), .S(n4291), .Z(
        n9479) );
  CMXI2X1 U19176 ( .A0(n9479), .A1(n9473), .S(n4012), .Z(n9486) );
  CMX2X1 U19177 ( .A0(n9474), .A1(n9486), .S(n3808), .Z(n9501) );
  CMXI2X1 U19178 ( .A0(n9475), .A1(n9501), .S(n3284), .Z(N3039) );
  CMX2X1 U19179 ( .A0(mem_data1[978]), .A1(mem_data1[979]), .S(n4291), .Z(
        n9482) );
  CMXI2X1 U19180 ( .A0(n9482), .A1(n9476), .S(n4011), .Z(n9489) );
  CMX2X1 U19181 ( .A0(n9477), .A1(n9489), .S(n3809), .Z(n9504) );
  CMXI2X1 U19182 ( .A0(n9478), .A1(n9504), .S(n3284), .Z(N3040) );
  CMX2X1 U19183 ( .A0(mem_data1[979]), .A1(mem_data1[980]), .S(n4291), .Z(
        n9485) );
  CMXI2X1 U19184 ( .A0(n9485), .A1(n9479), .S(n4011), .Z(n9492) );
  CMX2X1 U19185 ( .A0(n9480), .A1(n9492), .S(n3810), .Z(n9507) );
  CMXI2X1 U19186 ( .A0(n9481), .A1(n9507), .S(n3284), .Z(N3041) );
  CMX2X1 U19187 ( .A0(mem_data1[980]), .A1(mem_data1[981]), .S(n4290), .Z(
        n9488) );
  CMXI2X1 U19188 ( .A0(n9488), .A1(n9482), .S(n4011), .Z(n9497) );
  CMX2X1 U19189 ( .A0(n9483), .A1(n9497), .S(n3811), .Z(n9510) );
  CMXI2X1 U19190 ( .A0(n9484), .A1(n9510), .S(n3285), .Z(N3042) );
  CMX2X1 U19191 ( .A0(mem_data1[981]), .A1(mem_data1[982]), .S(n4290), .Z(
        n9491) );
  CMXI2X1 U19192 ( .A0(n9491), .A1(n9485), .S(n4011), .Z(n9500) );
  CMX2X1 U19193 ( .A0(n9486), .A1(n9500), .S(n3812), .Z(n9513) );
  CMXI2X1 U19194 ( .A0(n9487), .A1(n9513), .S(n3285), .Z(N3043) );
  CMX2X1 U19195 ( .A0(mem_data1[982]), .A1(mem_data1[983]), .S(n4290), .Z(
        n9496) );
  CMXI2X1 U19196 ( .A0(n9496), .A1(n9488), .S(n4011), .Z(n9503) );
  CMX2X1 U19197 ( .A0(n9489), .A1(n9503), .S(n4353), .Z(n9516) );
  CMXI2X1 U19198 ( .A0(n9490), .A1(n9516), .S(n3285), .Z(N3044) );
  CMX2X1 U19199 ( .A0(mem_data1[983]), .A1(mem_data1[984]), .S(n4290), .Z(
        n9499) );
  CMXI2X1 U19200 ( .A0(n9499), .A1(n9491), .S(n4011), .Z(n9506) );
  CMX2X1 U19201 ( .A0(n9492), .A1(n9506), .S(n3771), .Z(n9519) );
  CMXI2X1 U19202 ( .A0(n9493), .A1(n9519), .S(n3285), .Z(N3045) );
  CMXI2X1 U19203 ( .A0(n9495), .A1(n9494), .S(n3282), .Z(N2172) );
  CMX2X1 U19204 ( .A0(mem_data1[984]), .A1(mem_data1[985]), .S(n4290), .Z(
        n9502) );
  CMXI2X1 U19205 ( .A0(n9502), .A1(n9496), .S(n4011), .Z(n9509) );
  CMX2X1 U19206 ( .A0(n9497), .A1(n9509), .S(n3776), .Z(n9522) );
  CMXI2X1 U19207 ( .A0(n9498), .A1(n9522), .S(n3282), .Z(N3046) );
  CMX2X1 U19208 ( .A0(mem_data1[985]), .A1(mem_data1[986]), .S(n4290), .Z(
        n9505) );
  CMXI2X1 U19209 ( .A0(n9505), .A1(n9499), .S(n4011), .Z(n9512) );
  CMX2X1 U19210 ( .A0(n9500), .A1(n9512), .S(n3775), .Z(n9525) );
  CMXI2X1 U19211 ( .A0(n9501), .A1(n9525), .S(n3282), .Z(N3047) );
  CMX2X1 U19212 ( .A0(mem_data1[986]), .A1(mem_data1[987]), .S(n4290), .Z(
        n9508) );
  CMXI2X1 U19213 ( .A0(n9508), .A1(n9502), .S(n4011), .Z(n9515) );
  CMX2X1 U19214 ( .A0(n9503), .A1(n9515), .S(n3808), .Z(n9530) );
  CMXI2X1 U19215 ( .A0(n9504), .A1(n9530), .S(n3282), .Z(N3048) );
  CMX2X1 U19216 ( .A0(mem_data1[987]), .A1(mem_data1[988]), .S(n4290), .Z(
        n9511) );
  CMXI2X1 U19217 ( .A0(n9511), .A1(n9505), .S(n4011), .Z(n9518) );
  CMX2X1 U19218 ( .A0(n9506), .A1(n9518), .S(n3809), .Z(n9533) );
  CMXI2X1 U19219 ( .A0(n9507), .A1(n9533), .S(n3282), .Z(N3049) );
  CMX2X1 U19220 ( .A0(mem_data1[988]), .A1(mem_data1[989]), .S(n4290), .Z(
        n9514) );
  CMXI2X1 U19221 ( .A0(n9514), .A1(n9508), .S(n4011), .Z(n9521) );
  CMX2X1 U19222 ( .A0(n9509), .A1(n9521), .S(n3810), .Z(n9536) );
  CMXI2X1 U19223 ( .A0(n9510), .A1(n9536), .S(n3282), .Z(N3050) );
  CMX2X1 U19224 ( .A0(mem_data1[989]), .A1(mem_data1[990]), .S(n4290), .Z(
        n9517) );
  CMXI2X1 U19225 ( .A0(n9517), .A1(n9511), .S(n4011), .Z(n9524) );
  CMX2X1 U19226 ( .A0(n9512), .A1(n9524), .S(n3811), .Z(n9539) );
  CMXI2X1 U19227 ( .A0(n9513), .A1(n9539), .S(n3282), .Z(N3051) );
  CMX2X1 U19228 ( .A0(mem_data1[990]), .A1(mem_data1[991]), .S(n4290), .Z(
        n9520) );
  CMXI2X1 U19229 ( .A0(n9520), .A1(n9514), .S(n4011), .Z(n9529) );
  CMX2X1 U19230 ( .A0(n9515), .A1(n9529), .S(n3812), .Z(n9542) );
  CMXI2X1 U19231 ( .A0(n9516), .A1(n9542), .S(n3282), .Z(N3052) );
  CMX2X1 U19232 ( .A0(mem_data1[991]), .A1(mem_data1[992]), .S(n4289), .Z(
        n9523) );
  CMXI2X1 U19233 ( .A0(n9523), .A1(n9517), .S(n4011), .Z(n9532) );
  CMX2X1 U19234 ( .A0(n9518), .A1(n9532), .S(n3806), .Z(n9545) );
  CMXI2X1 U19235 ( .A0(n9519), .A1(n9545), .S(n3282), .Z(N3053) );
  CMX2X1 U19236 ( .A0(mem_data1[992]), .A1(mem_data1[993]), .S(n4289), .Z(
        n9528) );
  CMXI2X1 U19237 ( .A0(n9528), .A1(n9520), .S(n4011), .Z(n9535) );
  CMX2X1 U19238 ( .A0(n9521), .A1(n9535), .S(n3772), .Z(n9549) );
  CMXI2X1 U19239 ( .A0(n9522), .A1(n9549), .S(n3282), .Z(N3054) );
  CMX2X1 U19240 ( .A0(mem_data1[993]), .A1(mem_data1[994]), .S(n4289), .Z(
        n9531) );
  CMXI2X1 U19241 ( .A0(n9531), .A1(n9523), .S(n4011), .Z(n9538) );
  CMX2X1 U19242 ( .A0(n9524), .A1(n9538), .S(n3773), .Z(n9553) );
  CMXI2X1 U19243 ( .A0(n9525), .A1(n9553), .S(n3283), .Z(N3055) );
  CMXI2X1 U19244 ( .A0(n9527), .A1(n9526), .S(n3283), .Z(N2173) );
  CMX2X1 U19245 ( .A0(mem_data1[994]), .A1(mem_data1[995]), .S(n4289), .Z(
        n9534) );
  CMXI2X1 U19246 ( .A0(n9534), .A1(n9528), .S(n4010), .Z(n9541) );
  CMX2X1 U19247 ( .A0(n9529), .A1(n9541), .S(n3774), .Z(n9556) );
  CMXI2X1 U19248 ( .A0(n9530), .A1(n9556), .S(n3283), .Z(N3056) );
  CMX2X1 U19249 ( .A0(mem_data1[995]), .A1(mem_data1[996]), .S(n4289), .Z(
        n9537) );
  CMXI2X1 U19250 ( .A0(n9537), .A1(n9531), .S(n4010), .Z(n9544) );
  CMX2X1 U19251 ( .A0(n9532), .A1(n9544), .S(n3775), .Z(n9559) );
  CMXI2X1 U19252 ( .A0(n9533), .A1(n9559), .S(n3283), .Z(N3057) );
  CMX2X1 U19253 ( .A0(mem_data1[996]), .A1(mem_data1[997]), .S(n4289), .Z(
        n9540) );
  CMXI2X1 U19254 ( .A0(n9540), .A1(n9534), .S(n4010), .Z(n9548) );
  CMX2X1 U19255 ( .A0(n9535), .A1(n9548), .S(n3776), .Z(n9564) );
  CMXI2X1 U19256 ( .A0(n9536), .A1(n9564), .S(n3283), .Z(N3058) );
  CMX2X1 U19257 ( .A0(mem_data1[997]), .A1(mem_data1[998]), .S(n4289), .Z(
        n9543) );
  CMXI2X1 U19258 ( .A0(n9543), .A1(n9537), .S(n4010), .Z(n9552) );
  CMX2X1 U19259 ( .A0(n9538), .A1(n9552), .S(n3777), .Z(n9567) );
  CMXI2X1 U19260 ( .A0(n9539), .A1(n9567), .S(n3283), .Z(N3059) );
  CMX2X1 U19261 ( .A0(mem_data1[998]), .A1(mem_data1[999]), .S(n4289), .Z(
        n9546) );
  CMXI2X1 U19262 ( .A0(n9546), .A1(n9540), .S(n4010), .Z(n9555) );
  CMX2X1 U19263 ( .A0(n9541), .A1(n9555), .S(n3790), .Z(n9569) );
  CMXI2X1 U19264 ( .A0(n9542), .A1(n9569), .S(n3283), .Z(N3060) );
  CMX2X1 U19265 ( .A0(mem_data1[999]), .A1(mem_data1[1000]), .S(n4289), .Z(
        n9550) );
  CMXI2X1 U19266 ( .A0(n9550), .A1(n9543), .S(n4010), .Z(n9558) );
  CMX2X1 U19267 ( .A0(n9544), .A1(n9558), .S(n3791), .Z(n9571) );
  CMXI2X1 U19268 ( .A0(n9545), .A1(n9571), .S(n3280), .Z(N3061) );
  CMXI2X1 U19269 ( .A0(n9547), .A1(n9546), .S(n4010), .Z(n9563) );
  CMX2X1 U19270 ( .A0(n9548), .A1(n9563), .S(n3792), .Z(n9573) );
  CMXI2X1 U19271 ( .A0(n9549), .A1(n9573), .S(n3280), .Z(N3062) );
  CMXI2X1 U19272 ( .A0(n9551), .A1(n9550), .S(n4010), .Z(n9566) );
  CMX2X1 U19273 ( .A0(n9552), .A1(n9566), .S(n3793), .Z(n9575) );
  CMXI2X1 U19274 ( .A0(n9553), .A1(n9575), .S(n3280), .Z(N3063) );
  CMX2X1 U19275 ( .A0(n9555), .A1(n9554), .S(n3794), .Z(n9577) );
  CMXI2X1 U19276 ( .A0(n9556), .A1(n9577), .S(n3280), .Z(N3064) );
  CMX2X1 U19277 ( .A0(n9558), .A1(n9557), .S(n3795), .Z(n9579) );
  CMXI2X1 U19278 ( .A0(n9559), .A1(n9579), .S(n3280), .Z(N3065) );
  CMXI2X1 U19279 ( .A0(n9561), .A1(n9560), .S(n3280), .Z(N2174) );
  CMX2X1 U19280 ( .A0(n9563), .A1(n9562), .S(n3796), .Z(n9581) );
  CMXI2X1 U19281 ( .A0(n9564), .A1(n9581), .S(n3281), .Z(N3066) );
  CMX2X1 U19282 ( .A0(n9566), .A1(n9565), .S(n3797), .Z(n9583) );
  CMXI2X1 U19283 ( .A0(n9567), .A1(n9583), .S(n3281), .Z(N3067) );
  CMXI2X1 U19284 ( .A0(n9569), .A1(n9568), .S(n3281), .Z(N3068) );
  CMXI2X1 U19285 ( .A0(n9571), .A1(n9570), .S(n3281), .Z(N3069) );
  CMXI2X1 U19286 ( .A0(n9573), .A1(n9572), .S(n3281), .Z(N3070) );
  CMXI2X1 U19287 ( .A0(n9575), .A1(n9574), .S(n3281), .Z(N3071) );
  CMXI2X1 U19288 ( .A0(n9577), .A1(n9576), .S(n3281), .Z(N3072) );
  CMXI2X1 U19289 ( .A0(n9579), .A1(n9578), .S(n3281), .Z(N3073) );
  CMXI2X1 U19290 ( .A0(n9581), .A1(n9580), .S(n3281), .Z(N3074) );
  CMXI2X1 U19291 ( .A0(n9583), .A1(n9582), .S(n3281), .Z(N3075) );
  CMXI2X1 U19292 ( .A0(n9585), .A1(n9584), .S(n3281), .Z(N2175) );
  CMXI2X1 U19293 ( .A0(n9587), .A1(n9586), .S(n3282), .Z(N2085) );
  CMXI2X1 U19294 ( .A0(N8272), .A1(N8273), .S(n3884), .Z(n10328) );
  CMXI2X1 U19295 ( .A0(N8274), .A1(N8275), .S(n3886), .Z(n10331) );
  CMXI2X1 U19296 ( .A0(n10328), .A1(n10331), .S(n4138), .Z(n11003) );
  CMXI2X1 U19297 ( .A0(N8277), .A1(N8276), .S(n3869), .Z(n10330) );
  CMXI2X1 U19298 ( .A0(N8278), .A1(N8279), .S(n3888), .Z(n9588) );
  CMXI2X1 U19299 ( .A0(n10330), .A1(n9588), .S(n4138), .Z(n9589) );
  CMXI2X1 U19300 ( .A0(n11003), .A1(n9589), .S(n3801), .Z(n9590) );
  CMX2X1 U19301 ( .A0(N8269), .A1(N8268), .S(n4289), .Z(n9685) );
  CMXI2X1 U19302 ( .A0(N8270), .A1(N8271), .S(n3888), .Z(n10329) );
  CMXI2X1 U19303 ( .A0(n9685), .A1(n4432), .S(n4138), .Z(n11002) );
  CMX2X1 U19304 ( .A0(N8265), .A1(N8264), .S(n4289), .Z(n9687) );
  CMX2X1 U19305 ( .A0(N8267), .A1(N8266), .S(n4288), .Z(n9686) );
  CMXI2X1 U19306 ( .A0(n9687), .A1(n9686), .S(n4138), .Z(n9750) );
  CMX2X1 U19307 ( .A0(n11002), .A1(n9750), .S(n3791), .Z(n12341) );
  CMXI2X1 U19308 ( .A0(n9590), .A1(n12341), .S(n3499), .Z(N5158) );
  CMX2X1 U19309 ( .A0(N7277), .A1(N7276), .S(n4288), .Z(n9591) );
  CMXI2X1 U19310 ( .A0(n9591), .A1(n12619), .S(n4137), .Z(n12626) );
  CMX2X1 U19311 ( .A0(N7275), .A1(N7274), .S(n4288), .Z(n9592) );
  CMXI2X1 U19312 ( .A0(n9593), .A1(n9592), .S(n4137), .Z(n9606) );
  CMX2X1 U19313 ( .A0(n12626), .A1(n9606), .S(n3772), .Z(n12640) );
  CMXI2X1 U19314 ( .A0(n9595), .A1(n9594), .S(n4137), .Z(n9605) );
  CMXI2X1 U19315 ( .A0(n9597), .A1(n9596), .S(n4137), .Z(n9608) );
  CMX2X1 U19316 ( .A0(n9605), .A1(n9608), .S(n3773), .Z(n9623) );
  CMXI2X1 U19317 ( .A0(n12640), .A1(n9623), .S(n3499), .Z(N6158) );
  CMX2X1 U19318 ( .A0(N7276), .A1(N7275), .S(n4288), .Z(n9598) );
  CMX2X1 U19319 ( .A0(N7278), .A1(N7277), .S(n4288), .Z(n12623) );
  CMXI2X1 U19320 ( .A0(n9598), .A1(n12623), .S(n4137), .Z(n12629) );
  CMX2X1 U19321 ( .A0(N7274), .A1(N7273), .S(n4287), .Z(n9599) );
  CMXI2X1 U19322 ( .A0(n9600), .A1(n9599), .S(n4137), .Z(n9610) );
  CMX2X1 U19323 ( .A0(n12629), .A1(n9610), .S(n3774), .Z(n12642) );
  CMXI2X1 U19324 ( .A0(n9602), .A1(n9601), .S(n4137), .Z(n9609) );
  CMXI2X1 U19325 ( .A0(n9604), .A1(n9603), .S(n4137), .Z(n9612) );
  CMX2X1 U19326 ( .A0(n9609), .A1(n9612), .S(n3775), .Z(n9626) );
  CMXI2X1 U19327 ( .A0(n12642), .A1(n9626), .S(n3500), .Z(N6159) );
  CMXI2X1 U19328 ( .A0(n9592), .A1(n9591), .S(n4137), .Z(n12634) );
  CMXI2X1 U19329 ( .A0(n9594), .A1(n9593), .S(n4137), .Z(n9614) );
  CMX2X1 U19330 ( .A0(n12634), .A1(n9614), .S(n3776), .Z(n12644) );
  CMXI2X1 U19331 ( .A0(n9596), .A1(n9595), .S(n4137), .Z(n9613) );
  CMXI2X1 U19332 ( .A0(n9607), .A1(n9597), .S(n4137), .Z(n9616) );
  CMX2X1 U19333 ( .A0(n9613), .A1(n9616), .S(n3777), .Z(n9629) );
  CMXI2X1 U19334 ( .A0(n12644), .A1(n9629), .S(n3500), .Z(N6160) );
  CMXI2X1 U19335 ( .A0(n9599), .A1(n9598), .S(n4137), .Z(n12637) );
  CMXI2X1 U19336 ( .A0(n9601), .A1(n9600), .S(n4137), .Z(n9618) );
  CMX2X1 U19337 ( .A0(n12637), .A1(n9618), .S(n3790), .Z(n12646) );
  CMXI2X1 U19338 ( .A0(n9603), .A1(n9602), .S(n4137), .Z(n9617) );
  CMXI2X1 U19339 ( .A0(n9611), .A1(n9604), .S(n4137), .Z(n9620) );
  CMX2X1 U19340 ( .A0(n9617), .A1(n9620), .S(n3791), .Z(n9632) );
  CMXI2X1 U19341 ( .A0(n12646), .A1(n9632), .S(n3500), .Z(N6161) );
  CMX2X1 U19342 ( .A0(n9606), .A1(n9605), .S(n3792), .Z(n12648) );
  CMXI2X1 U19343 ( .A0(n9615), .A1(n9607), .S(n4136), .Z(n9622) );
  CMX2X1 U19344 ( .A0(n9608), .A1(n9622), .S(n3793), .Z(n9634) );
  CMXI2X1 U19345 ( .A0(n12648), .A1(n9634), .S(n3500), .Z(N6162) );
  CMX2X1 U19346 ( .A0(n9610), .A1(n9609), .S(n3794), .Z(n12650) );
  CMXI2X1 U19347 ( .A0(n9619), .A1(n9611), .S(n4136), .Z(n9625) );
  CMX2X1 U19348 ( .A0(n9612), .A1(n9625), .S(n3795), .Z(n9636) );
  CMXI2X1 U19349 ( .A0(n12650), .A1(n9636), .S(n3500), .Z(N6163) );
  CMX2X1 U19350 ( .A0(n9614), .A1(n9613), .S(n3796), .Z(n12652) );
  CMXI2X1 U19351 ( .A0(n9621), .A1(n9615), .S(n4136), .Z(n9628) );
  CMX2X1 U19352 ( .A0(n9616), .A1(n9628), .S(n3797), .Z(n9638) );
  CMX2X1 U19353 ( .A0(n9618), .A1(n9617), .S(n3805), .Z(n12654) );
  CMXI2X1 U19354 ( .A0(n9624), .A1(n9619), .S(n4136), .Z(n9631) );
  CMX2X1 U19355 ( .A0(n9620), .A1(n9631), .S(n3806), .Z(n9640) );
  CMXI2X1 U19356 ( .A0(n12654), .A1(n9640), .S(n3500), .Z(N6165) );
  CMXI2X1 U19357 ( .A0(n9627), .A1(n9621), .S(n4136), .Z(n9633) );
  CMX2X1 U19358 ( .A0(n9622), .A1(n9633), .S(n3773), .Z(n9641) );
  CMXI2X1 U19359 ( .A0(n9623), .A1(n9641), .S(n3500), .Z(N6166) );
  CMXI2X1 U19360 ( .A0(n9630), .A1(n9624), .S(n4136), .Z(n9635) );
  CMX2X1 U19361 ( .A0(n9625), .A1(n9635), .S(n3774), .Z(n9642) );
  CMXI2X1 U19362 ( .A0(n9626), .A1(n9642), .S(n3500), .Z(N6167) );
  CMXI2X1 U19363 ( .A0(n9649), .A1(n12237), .S(n4136), .Z(n12304) );
  CMX2X1 U19364 ( .A0(N8173), .A1(N8172), .S(n4283), .Z(n9651) );
  CMXI2X1 U19365 ( .A0(n9651), .A1(n9650), .S(n4136), .Z(n9664) );
  CMX2X1 U19366 ( .A0(n12304), .A1(n9664), .S(n3809), .Z(n12438) );
  CMXI2X1 U19367 ( .A0(n9653), .A1(n9652), .S(n4136), .Z(n9663) );
  CMX2X1 U19368 ( .A0(N8167), .A1(N8166), .S(n4282), .Z(n9654) );
  CMXI2X1 U19369 ( .A0(n9655), .A1(n9654), .S(n4136), .Z(n9666) );
  CMX2X1 U19370 ( .A0(n9663), .A1(n9666), .S(n3810), .Z(n9681) );
  CMXI2X1 U19371 ( .A0(n12438), .A1(n9681), .S(n3500), .Z(N5258) );
  CMX2X1 U19372 ( .A0(n9628), .A1(n9637), .S(n3775), .Z(n9643) );
  CMXI2X1 U19373 ( .A0(n9629), .A1(n9643), .S(n3500), .Z(N6168) );
  CMX2X1 U19374 ( .A0(n9631), .A1(n9639), .S(n3776), .Z(n9644) );
  CMXI2X1 U19375 ( .A0(n9632), .A1(n9644), .S(n3501), .Z(N6169) );
  CMXI2X1 U19376 ( .A0(n9634), .A1(n9645), .S(n3501), .Z(N6170) );
  CMXI2X1 U19377 ( .A0(n9636), .A1(n9646), .S(n3501), .Z(N6171) );
  CMXI2X1 U19378 ( .A0(n9638), .A1(n9647), .S(n3501), .Z(N6172) );
  CND2IX1 U19379 ( .B(n9639), .A(n3802), .Z(n9648) );
  CMXI2X1 U19380 ( .A0(n9640), .A1(n9648), .S(n3499), .Z(N6173) );
  CMXI2X1 U19381 ( .A0(n9656), .A1(n12271), .S(n4136), .Z(n12337) );
  CMX2X1 U19382 ( .A0(N8172), .A1(N8171), .S(n4286), .Z(n9658) );
  CMX2X1 U19383 ( .A0(N8174), .A1(N8173), .S(n4286), .Z(n9657) );
  CMXI2X1 U19384 ( .A0(n9658), .A1(n9657), .S(n4136), .Z(n9668) );
  CMX2X1 U19385 ( .A0(n12337), .A1(n9668), .S(n3797), .Z(n12470) );
  CMX2X1 U19386 ( .A0(N8168), .A1(N8167), .S(n4286), .Z(n9660) );
  CMXI2X1 U19387 ( .A0(n9660), .A1(n9659), .S(n4136), .Z(n9667) );
  CMX2X1 U19388 ( .A0(N8166), .A1(N8165), .S(n4286), .Z(n9661) );
  CMXI2X1 U19389 ( .A0(n9662), .A1(n9661), .S(n4136), .Z(n9670) );
  CMX2X1 U19390 ( .A0(n9667), .A1(n9670), .S(n3805), .Z(n9684) );
  CMXI2X1 U19391 ( .A0(n12470), .A1(n9684), .S(n3501), .Z(N5259) );
  CMXI2X1 U19392 ( .A0(n9650), .A1(n9649), .S(n4136), .Z(n12372) );
  CMXI2X1 U19393 ( .A0(n9652), .A1(n9651), .S(n4136), .Z(n9672) );
  CMX2X1 U19394 ( .A0(n12372), .A1(n9672), .S(n3806), .Z(n12502) );
  CMXI2X1 U19395 ( .A0(n9654), .A1(n9653), .S(n4135), .Z(n9671) );
  CMXI2X1 U19396 ( .A0(n9665), .A1(n9655), .S(n4135), .Z(n9674) );
  CMX2X1 U19397 ( .A0(n9671), .A1(n9674), .S(n3807), .Z(n9690) );
  CMXI2X1 U19398 ( .A0(n12502), .A1(n9690), .S(n3499), .Z(N5260) );
  CMXI2X1 U19399 ( .A0(n9657), .A1(n9656), .S(n4135), .Z(n12405) );
  CMXI2X1 U19400 ( .A0(n9659), .A1(n9658), .S(n4135), .Z(n9676) );
  CMX2X1 U19401 ( .A0(n12405), .A1(n9676), .S(n3808), .Z(n12534) );
  CMXI2X1 U19402 ( .A0(n9661), .A1(n9660), .S(n4135), .Z(n9675) );
  CMXI2X1 U19403 ( .A0(n9669), .A1(n9662), .S(n4135), .Z(n9678) );
  CMX2X1 U19404 ( .A0(n9675), .A1(n9678), .S(n3792), .Z(n9693) );
  CMXI2X1 U19405 ( .A0(n12534), .A1(n9693), .S(n3499), .Z(N5261) );
  CMX2X1 U19406 ( .A0(n9664), .A1(n9663), .S(n3807), .Z(n12566) );
  CMXI2X1 U19407 ( .A0(n9673), .A1(n9665), .S(n4135), .Z(n9680) );
  CMX2X1 U19408 ( .A0(n9666), .A1(n9680), .S(n3808), .Z(n9696) );
  CMXI2X1 U19409 ( .A0(n12566), .A1(n9696), .S(n3499), .Z(N5262) );
  CMX2X1 U19410 ( .A0(n9668), .A1(n9667), .S(n3810), .Z(n12598) );
  CMX2X1 U19411 ( .A0(N8160), .A1(N8159), .S(n4285), .Z(n9677) );
  CMXI2X1 U19412 ( .A0(n9677), .A1(n9669), .S(n4135), .Z(n9683) );
  CMX2X1 U19413 ( .A0(n9670), .A1(n9683), .S(n3811), .Z(n9699) );
  CMXI2X1 U19414 ( .A0(n12598), .A1(n9699), .S(n3499), .Z(N5263) );
  CMX2X1 U19415 ( .A0(n9672), .A1(n9671), .S(n3812), .Z(n12632) );
  CMXI2X1 U19416 ( .A0(n9679), .A1(n9673), .S(n4135), .Z(n9689) );
  CMX2X1 U19417 ( .A0(n9674), .A1(n9689), .S(n4324), .Z(n9702) );
  CMXI2X1 U19418 ( .A0(n12632), .A1(n9702), .S(n3283), .Z(N5264) );
  CMX2X1 U19419 ( .A0(n9676), .A1(n9675), .S(n3771), .Z(n12656) );
  CMXI2X1 U19420 ( .A0(n9682), .A1(n9677), .S(n4135), .Z(n9692) );
  CMX2X1 U19421 ( .A0(n9678), .A1(n9692), .S(n3772), .Z(n9705) );
  CMXI2X1 U19422 ( .A0(n12656), .A1(n9705), .S(n3285), .Z(N5265) );
  CMXI2X1 U19423 ( .A0(n9688), .A1(n9679), .S(n4135), .Z(n9695) );
  CMX2X1 U19424 ( .A0(n9680), .A1(n9695), .S(n3773), .Z(n9708) );
  CMXI2X1 U19425 ( .A0(n9681), .A1(n9708), .S(n3503), .Z(N5266) );
  CMXI2X1 U19426 ( .A0(n9691), .A1(n9682), .S(n4135), .Z(n9698) );
  CMX2X1 U19427 ( .A0(n9683), .A1(n9698), .S(n3774), .Z(n9711) );
  CMXI2X1 U19428 ( .A0(n9684), .A1(n9711), .S(n3502), .Z(N5267) );
  CMXI2X1 U19429 ( .A0(n9686), .A1(n9685), .S(n4135), .Z(n11670) );
  CMX2X1 U19430 ( .A0(N8263), .A1(N8262), .S(n4285), .Z(n9748) );
  CMXI2X1 U19431 ( .A0(n9748), .A1(n9687), .S(n4135), .Z(n9822) );
  CMX2X1 U19432 ( .A0(n11670), .A1(n9822), .S(n3775), .Z(n10333) );
  CMX2X1 U19433 ( .A0(N8259), .A1(N8258), .S(n4285), .Z(n9751) );
  CMX2X1 U19434 ( .A0(N8261), .A1(N8260), .S(n4285), .Z(n9749) );
  CMXI2X1 U19435 ( .A0(n9751), .A1(n9749), .S(n4135), .Z(n9821) );
  CMX2X1 U19436 ( .A0(N8255), .A1(N8254), .S(n4285), .Z(n9753) );
  CMX2X1 U19437 ( .A0(N8257), .A1(N8256), .S(n4285), .Z(n9752) );
  CMXI2X1 U19438 ( .A0(n9753), .A1(n9752), .S(n4135), .Z(n9824) );
  CMX2X1 U19439 ( .A0(n9821), .A1(n9824), .S(n3776), .Z(n9959) );
  CMXI2X1 U19440 ( .A0(n10333), .A1(n9959), .S(n3502), .Z(N5168) );
  CMXI2X1 U19441 ( .A0(n9694), .A1(n9688), .S(n4134), .Z(n9701) );
  CMX2X1 U19442 ( .A0(n9689), .A1(n9701), .S(n3777), .Z(n9714) );
  CMXI2X1 U19443 ( .A0(n9690), .A1(n9714), .S(n3502), .Z(N5268) );
  CMXI2X1 U19444 ( .A0(n9697), .A1(n9691), .S(n4134), .Z(n9704) );
  CMX2X1 U19445 ( .A0(n9692), .A1(n9704), .S(n3790), .Z(n9717) );
  CMXI2X1 U19446 ( .A0(n9693), .A1(n9717), .S(n3502), .Z(N5269) );
  CMXI2X1 U19447 ( .A0(n9700), .A1(n9694), .S(n4134), .Z(n9707) );
  CMX2X1 U19448 ( .A0(n9695), .A1(n9707), .S(n3791), .Z(n9720) );
  CMXI2X1 U19449 ( .A0(n9696), .A1(n9720), .S(n3502), .Z(N5270) );
  CMXI2X1 U19450 ( .A0(n9703), .A1(n9697), .S(n4134), .Z(n9710) );
  CMX2X1 U19451 ( .A0(n9698), .A1(n9710), .S(n3810), .Z(n9723) );
  CMXI2X1 U19452 ( .A0(n9699), .A1(n9723), .S(n3502), .Z(N5271) );
  CMX2X1 U19453 ( .A0(N8151), .A1(N8150), .S(n4284), .Z(n9706) );
  CMXI2X1 U19454 ( .A0(n9706), .A1(n9700), .S(n4134), .Z(n9713) );
  CMX2X1 U19455 ( .A0(n9701), .A1(n9713), .S(n3811), .Z(n9726) );
  CMXI2X1 U19456 ( .A0(n9702), .A1(n9726), .S(n3502), .Z(N5272) );
  CMX2X1 U19457 ( .A0(N8150), .A1(N8149), .S(n4284), .Z(n9709) );
  CMXI2X1 U19458 ( .A0(n9709), .A1(n9703), .S(n4134), .Z(n9716) );
  CMX2X1 U19459 ( .A0(n9704), .A1(n9716), .S(n3809), .Z(n9729) );
  CMXI2X1 U19460 ( .A0(n9705), .A1(n9729), .S(n3502), .Z(N5273) );
  CMX2X1 U19461 ( .A0(N8149), .A1(N8148), .S(n4284), .Z(n9712) );
  CMXI2X1 U19462 ( .A0(n9712), .A1(n9706), .S(n4134), .Z(n9719) );
  CMX2X1 U19463 ( .A0(n9707), .A1(n9719), .S(n3810), .Z(n9732) );
  CMXI2X1 U19464 ( .A0(n9708), .A1(n9732), .S(n3502), .Z(N5274) );
  CMX2X1 U19465 ( .A0(N8148), .A1(N8147), .S(n4284), .Z(n9715) );
  CMXI2X1 U19466 ( .A0(n9715), .A1(n9709), .S(n4134), .Z(n9722) );
  CMX2X1 U19467 ( .A0(n9710), .A1(n9722), .S(n3811), .Z(n9735) );
  CMXI2X1 U19468 ( .A0(n9711), .A1(n9735), .S(n3502), .Z(N5275) );
  CMX2X1 U19469 ( .A0(N8147), .A1(N8146), .S(n4284), .Z(n9718) );
  CMXI2X1 U19470 ( .A0(n9718), .A1(n9712), .S(n4134), .Z(n9725) );
  CMX2X1 U19471 ( .A0(n9713), .A1(n9725), .S(n3812), .Z(n9738) );
  CMXI2X1 U19472 ( .A0(n9714), .A1(n9738), .S(n3502), .Z(N5276) );
  CMX2X1 U19473 ( .A0(N8146), .A1(N8145), .S(n4284), .Z(n9721) );
  CMXI2X1 U19474 ( .A0(n9721), .A1(n9715), .S(n4134), .Z(n9728) );
  CMX2X1 U19475 ( .A0(n9716), .A1(n9728), .S(n4316), .Z(n9741) );
  CMXI2X1 U19476 ( .A0(n9717), .A1(n9741), .S(n3501), .Z(N5277) );
  CMX2X1 U19477 ( .A0(N8266), .A1(N8265), .S(n4284), .Z(n9784) );
  CMX2X1 U19478 ( .A0(N8268), .A1(N8267), .S(n4284), .Z(n9995) );
  CMXI2X1 U19479 ( .A0(n9784), .A1(n9995), .S(n4134), .Z(n12004) );
  CMX2X1 U19480 ( .A0(N8262), .A1(N8261), .S(n4283), .Z(n9786) );
  CMX2X1 U19481 ( .A0(N8264), .A1(N8263), .S(n4283), .Z(n9785) );
  CMXI2X1 U19482 ( .A0(n9786), .A1(n9785), .S(n4134), .Z(n9856) );
  CMX2X1 U19483 ( .A0(n12004), .A1(n9856), .S(n3793), .Z(n10670) );
  CMX2X1 U19484 ( .A0(N8258), .A1(N8257), .S(n4283), .Z(n9788) );
  CMX2X1 U19485 ( .A0(N8260), .A1(N8259), .S(n4283), .Z(n9787) );
  CMXI2X1 U19486 ( .A0(n9788), .A1(n9787), .S(n4134), .Z(n9855) );
  CMX2X1 U19487 ( .A0(N8254), .A1(N8253), .S(n4283), .Z(n9790) );
  CMX2X1 U19488 ( .A0(N8256), .A1(N8255), .S(n4283), .Z(n9789) );
  CMXI2X1 U19489 ( .A0(n9790), .A1(n9789), .S(n4134), .Z(n9858) );
  CMX2X1 U19490 ( .A0(n9855), .A1(n9858), .S(n3792), .Z(n9992) );
  CMXI2X1 U19491 ( .A0(n10670), .A1(n9992), .S(n3501), .Z(N5169) );
  CMX2X1 U19492 ( .A0(N8145), .A1(N8144), .S(n4283), .Z(n9724) );
  CMXI2X1 U19493 ( .A0(n9724), .A1(n9718), .S(n4134), .Z(n9731) );
  CMX2X1 U19494 ( .A0(n9719), .A1(n9731), .S(n3793), .Z(n9744) );
  CMXI2X1 U19495 ( .A0(n9720), .A1(n9744), .S(n3501), .Z(N5278) );
  CMX2X1 U19496 ( .A0(N8144), .A1(N8143), .S(n4283), .Z(n9727) );
  CMXI2X1 U19497 ( .A0(n9727), .A1(n9721), .S(n4134), .Z(n9734) );
  CMX2X1 U19498 ( .A0(n9722), .A1(n9734), .S(n3794), .Z(n9747) );
  CMXI2X1 U19499 ( .A0(n9723), .A1(n9747), .S(n3501), .Z(N5279) );
  CMX2X1 U19500 ( .A0(N8143), .A1(N8142), .S(n4283), .Z(n9730) );
  CMXI2X1 U19501 ( .A0(n9730), .A1(n9724), .S(n4133), .Z(n9737) );
  CMX2X1 U19502 ( .A0(n9725), .A1(n9737), .S(n3795), .Z(n9756) );
  CMXI2X1 U19503 ( .A0(n9726), .A1(n9756), .S(n3501), .Z(N5280) );
  CMX2X1 U19504 ( .A0(N8142), .A1(N8141), .S(n4283), .Z(n9733) );
  CMXI2X1 U19505 ( .A0(n9733), .A1(n9727), .S(n4133), .Z(n9740) );
  CMX2X1 U19506 ( .A0(n9728), .A1(n9740), .S(n3796), .Z(n9759) );
  CMXI2X1 U19507 ( .A0(n9729), .A1(n9759), .S(n3501), .Z(N5281) );
  CMX2X1 U19508 ( .A0(N8141), .A1(N8140), .S(n4283), .Z(n9736) );
  CMXI2X1 U19509 ( .A0(n9736), .A1(n9730), .S(n4133), .Z(n9743) );
  CMX2X1 U19510 ( .A0(n9731), .A1(n9743), .S(n3797), .Z(n9762) );
  CMXI2X1 U19511 ( .A0(n9732), .A1(n9762), .S(n3504), .Z(N5282) );
  CMX2X1 U19512 ( .A0(N8140), .A1(N8139), .S(n4282), .Z(n9739) );
  CMXI2X1 U19513 ( .A0(n9739), .A1(n9733), .S(n4133), .Z(n9746) );
  CMX2X1 U19514 ( .A0(n9734), .A1(n9746), .S(n3805), .Z(n9765) );
  CMXI2X1 U19515 ( .A0(n9735), .A1(n9765), .S(n3504), .Z(N5283) );
  CMX2X1 U19516 ( .A0(N8139), .A1(N8138), .S(n4282), .Z(n9742) );
  CMXI2X1 U19517 ( .A0(n9742), .A1(n9736), .S(n4133), .Z(n9755) );
  CMX2X1 U19518 ( .A0(n9737), .A1(n9755), .S(n3806), .Z(n9768) );
  CMXI2X1 U19519 ( .A0(n9738), .A1(n9768), .S(n3504), .Z(N5284) );
  CMX2X1 U19520 ( .A0(N8138), .A1(N8137), .S(n4282), .Z(n9745) );
  CMXI2X1 U19521 ( .A0(n9745), .A1(n9739), .S(n4133), .Z(n9758) );
  CMX2X1 U19522 ( .A0(n9740), .A1(n9758), .S(n3807), .Z(n9771) );
  CMXI2X1 U19523 ( .A0(n9741), .A1(n9771), .S(n3504), .Z(N5285) );
  CMX2X1 U19524 ( .A0(N8137), .A1(N8136), .S(n4282), .Z(n9754) );
  CMXI2X1 U19525 ( .A0(n9754), .A1(n9742), .S(n4133), .Z(n9761) );
  CMX2X1 U19526 ( .A0(n9743), .A1(n9761), .S(n3808), .Z(n9774) );
  CMXI2X1 U19527 ( .A0(n9744), .A1(n9774), .S(n3504), .Z(N5286) );
  CMX2X1 U19528 ( .A0(N8136), .A1(N8135), .S(n4282), .Z(n9757) );
  CMXI2X1 U19529 ( .A0(n9757), .A1(n9745), .S(n4133), .Z(n9764) );
  CMX2X1 U19530 ( .A0(n9746), .A1(n9764), .S(n3809), .Z(n9777) );
  CMXI2X1 U19531 ( .A0(n9747), .A1(n9777), .S(n3504), .Z(N5287) );
  CMXI2X1 U19532 ( .A0(n9749), .A1(n9748), .S(n4133), .Z(n9890) );
  CMX2X1 U19533 ( .A0(n9750), .A1(n9890), .S(n3810), .Z(n11004) );
  CMXI2X1 U19534 ( .A0(n9752), .A1(n9751), .S(n4133), .Z(n9889) );
  CMX2X1 U19535 ( .A0(N8253), .A1(N8252), .S(n4282), .Z(n9823) );
  CMXI2X1 U19536 ( .A0(n9823), .A1(n9753), .S(n4133), .Z(n9892) );
  CMX2X1 U19537 ( .A0(n9889), .A1(n9892), .S(n3811), .Z(n10030) );
  CMXI2X1 U19538 ( .A0(n11004), .A1(n10030), .S(n3504), .Z(N5170) );
  CMX2X1 U19539 ( .A0(N8135), .A1(N8134), .S(n4282), .Z(n9760) );
  CMXI2X1 U19540 ( .A0(n9760), .A1(n9754), .S(n4133), .Z(n9767) );
  CMX2X1 U19541 ( .A0(n9755), .A1(n9767), .S(n3812), .Z(n9780) );
  CMXI2X1 U19542 ( .A0(n9756), .A1(n9780), .S(n3504), .Z(N5288) );
  CMX2X1 U19543 ( .A0(N8134), .A1(N8133), .S(n4282), .Z(n9763) );
  CMXI2X1 U19544 ( .A0(n9763), .A1(n9757), .S(n4133), .Z(n9770) );
  CMX2X1 U19545 ( .A0(n9758), .A1(n9770), .S(n4329), .Z(n9783) );
  CMXI2X1 U19546 ( .A0(n9759), .A1(n9783), .S(n3503), .Z(N5289) );
  CMX2X1 U19547 ( .A0(N8133), .A1(N8132), .S(n4282), .Z(n9766) );
  CMXI2X1 U19548 ( .A0(n9766), .A1(n9760), .S(n4133), .Z(n9773) );
  CMX2X1 U19549 ( .A0(n9761), .A1(n9773), .S(n3771), .Z(n9793) );
  CMXI2X1 U19550 ( .A0(n9762), .A1(n9793), .S(n3503), .Z(N5290) );
  CMX2X1 U19551 ( .A0(N8132), .A1(N8131), .S(n4282), .Z(n9769) );
  CMXI2X1 U19552 ( .A0(n9769), .A1(n9763), .S(n4133), .Z(n9776) );
  CMX2X1 U19553 ( .A0(n9764), .A1(n9776), .S(n3811), .Z(n9796) );
  CMXI2X1 U19554 ( .A0(n9765), .A1(n9796), .S(n3503), .Z(N5291) );
  CMX2X1 U19555 ( .A0(N8131), .A1(N8130), .S(n4282), .Z(n9772) );
  CMXI2X1 U19556 ( .A0(n9772), .A1(n9766), .S(n4133), .Z(n9779) );
  CMX2X1 U19557 ( .A0(n9767), .A1(n9779), .S(n3812), .Z(n9799) );
  CMXI2X1 U19558 ( .A0(n9768), .A1(n9799), .S(n3503), .Z(N5292) );
  CMX2X1 U19559 ( .A0(N8130), .A1(N8129), .S(n4281), .Z(n9775) );
  CMXI2X1 U19560 ( .A0(n9775), .A1(n9769), .S(n4132), .Z(n9782) );
  CMX2X1 U19561 ( .A0(n9770), .A1(n9782), .S(n3771), .Z(n9802) );
  CMXI2X1 U19562 ( .A0(n9771), .A1(n9802), .S(n3503), .Z(N5293) );
  CMX2X1 U19563 ( .A0(N8129), .A1(N8128), .S(n4281), .Z(n9778) );
  CMXI2X1 U19564 ( .A0(n9778), .A1(n9772), .S(n4132), .Z(n9792) );
  CMX2X1 U19565 ( .A0(n9773), .A1(n9792), .S(n3772), .Z(n9805) );
  CMXI2X1 U19566 ( .A0(n9774), .A1(n9805), .S(n3503), .Z(N5294) );
  CMX2X1 U19567 ( .A0(N8128), .A1(N8127), .S(n4281), .Z(n9781) );
  CMXI2X1 U19568 ( .A0(n9781), .A1(n9775), .S(n4132), .Z(n9795) );
  CMX2X1 U19569 ( .A0(n9776), .A1(n9795), .S(n3773), .Z(n9808) );
  CMXI2X1 U19570 ( .A0(n9777), .A1(n9808), .S(n3503), .Z(N5295) );
  CMX2X1 U19571 ( .A0(N8127), .A1(N8126), .S(n4281), .Z(n9791) );
  CMXI2X1 U19572 ( .A0(n9791), .A1(n9778), .S(n4132), .Z(n9798) );
  CMX2X1 U19573 ( .A0(n9779), .A1(n9798), .S(n3774), .Z(n9811) );
  CMXI2X1 U19574 ( .A0(n9780), .A1(n9811), .S(n3503), .Z(N5296) );
  CMX2X1 U19575 ( .A0(N8126), .A1(N8125), .S(n4281), .Z(n9794) );
  CMXI2X1 U19576 ( .A0(n9794), .A1(n9781), .S(n4132), .Z(n9801) );
  CMX2X1 U19577 ( .A0(n9782), .A1(n9801), .S(n3775), .Z(n9814) );
  CMXI2X1 U19578 ( .A0(n9783), .A1(n9814), .S(n3503), .Z(N5297) );
  CMXI2X1 U19579 ( .A0(n9785), .A1(n9784), .S(n4132), .Z(n9996) );
  CMXI2X1 U19580 ( .A0(n9787), .A1(n9786), .S(n4132), .Z(n9924) );
  CMX2X1 U19581 ( .A0(n9996), .A1(n9924), .S(n3794), .Z(n11338) );
  CMXI2X1 U19582 ( .A0(n9789), .A1(n9788), .S(n4132), .Z(n9923) );
  CMX2X1 U19583 ( .A0(N8252), .A1(N8251), .S(n4281), .Z(n9857) );
  CMXI2X1 U19584 ( .A0(n9857), .A1(n9790), .S(n4132), .Z(n9926) );
  CMX2X1 U19585 ( .A0(n9923), .A1(n9926), .S(n3772), .Z(n10063) );
  CMXI2X1 U19586 ( .A0(n11338), .A1(n10063), .S(n3503), .Z(N5171) );
  CMX2X1 U19587 ( .A0(N8125), .A1(N8124), .S(n4281), .Z(n9797) );
  CMXI2X1 U19588 ( .A0(n9797), .A1(n9791), .S(n4132), .Z(n9804) );
  CMX2X1 U19589 ( .A0(n9792), .A1(n9804), .S(n3773), .Z(n9817) );
  CMXI2X1 U19590 ( .A0(n9793), .A1(n9817), .S(n3506), .Z(N5298) );
  CMX2X1 U19591 ( .A0(N8124), .A1(N8123), .S(n4281), .Z(n9800) );
  CMXI2X1 U19592 ( .A0(n9800), .A1(n9794), .S(n4132), .Z(n9807) );
  CMX2X1 U19593 ( .A0(n9795), .A1(n9807), .S(n3774), .Z(n9820) );
  CMXI2X1 U19594 ( .A0(n9796), .A1(n9820), .S(n3506), .Z(N5299) );
  CMX2X1 U19595 ( .A0(N8123), .A1(N8122), .S(n4281), .Z(n9803) );
  CMXI2X1 U19596 ( .A0(n9803), .A1(n9797), .S(n4132), .Z(n9810) );
  CMX2X1 U19597 ( .A0(n9798), .A1(n9810), .S(n3775), .Z(n9827) );
  CMXI2X1 U19598 ( .A0(n9799), .A1(n9827), .S(n3506), .Z(N5300) );
  CMX2X1 U19599 ( .A0(N8122), .A1(N8121), .S(n4281), .Z(n9806) );
  CMXI2X1 U19600 ( .A0(n9806), .A1(n9800), .S(n4132), .Z(n9813) );
  CMX2X1 U19601 ( .A0(n9801), .A1(n9813), .S(n3809), .Z(n9830) );
  CMXI2X1 U19602 ( .A0(n9802), .A1(n9830), .S(n3506), .Z(N5301) );
  CMX2X1 U19603 ( .A0(N8121), .A1(N8120), .S(n4281), .Z(n9809) );
  CMXI2X1 U19604 ( .A0(n9809), .A1(n9803), .S(n4132), .Z(n9816) );
  CMX2X1 U19605 ( .A0(n9804), .A1(n9816), .S(n3808), .Z(n9833) );
  CMXI2X1 U19606 ( .A0(n9805), .A1(n9833), .S(n3505), .Z(N5302) );
  CMX2X1 U19607 ( .A0(N8120), .A1(N8119), .S(n4280), .Z(n9812) );
  CMXI2X1 U19608 ( .A0(n9812), .A1(n9806), .S(n4132), .Z(n9819) );
  CMX2X1 U19609 ( .A0(n9807), .A1(n9819), .S(n3809), .Z(n9836) );
  CMXI2X1 U19610 ( .A0(n9808), .A1(n9836), .S(n3505), .Z(N5303) );
  CMX2X1 U19611 ( .A0(N8119), .A1(N8118), .S(n4280), .Z(n9815) );
  CMXI2X1 U19612 ( .A0(n9815), .A1(n9809), .S(n4132), .Z(n9826) );
  CMX2X1 U19613 ( .A0(n9810), .A1(n9826), .S(n3810), .Z(n9839) );
  CMXI2X1 U19614 ( .A0(n9811), .A1(n9839), .S(n3505), .Z(N5304) );
  CMX2X1 U19615 ( .A0(N8118), .A1(N8117), .S(n4280), .Z(n9818) );
  CMXI2X1 U19616 ( .A0(n9818), .A1(n9812), .S(n4131), .Z(n9829) );
  CMX2X1 U19617 ( .A0(n9813), .A1(n9829), .S(n3811), .Z(n9842) );
  CMXI2X1 U19618 ( .A0(n9814), .A1(n9842), .S(n3505), .Z(N5305) );
  CMXI2X1 U19619 ( .A0(n9825), .A1(n9815), .S(n4131), .Z(n9832) );
  CMX2X1 U19620 ( .A0(n9816), .A1(n9832), .S(n3812), .Z(n9845) );
  CMXI2X1 U19621 ( .A0(n9817), .A1(n9845), .S(n3505), .Z(N5306) );
  CMXI2X1 U19622 ( .A0(n9828), .A1(n9818), .S(n4131), .Z(n9835) );
  CMX2X1 U19623 ( .A0(n9819), .A1(n9835), .S(n4311), .Z(n9848) );
  CMXI2X1 U19624 ( .A0(n9820), .A1(n9848), .S(n3505), .Z(N5307) );
  CMX2X1 U19625 ( .A0(n9822), .A1(n9821), .S(n3771), .Z(n11672) );
  CMX2X1 U19626 ( .A0(N8251), .A1(N8250), .S(n4280), .Z(n9891) );
  CMXI2X1 U19627 ( .A0(n9891), .A1(n9823), .S(n4131), .Z(n9958) );
  CMX2X1 U19628 ( .A0(n9824), .A1(n9958), .S(n3772), .Z(n10096) );
  CMXI2X1 U19629 ( .A0(n11672), .A1(n10096), .S(n3505), .Z(N5172) );
  CMX2X1 U19630 ( .A0(N8115), .A1(N8114), .S(n4280), .Z(n9831) );
  CMXI2X1 U19631 ( .A0(n9831), .A1(n9825), .S(n4131), .Z(n9838) );
  CMX2X1 U19632 ( .A0(n9826), .A1(n9838), .S(n3808), .Z(n9851) );
  CMXI2X1 U19633 ( .A0(n9827), .A1(n9851), .S(n3505), .Z(N5308) );
  CMX2X1 U19634 ( .A0(N8114), .A1(N8113), .S(n4280), .Z(n9834) );
  CMXI2X1 U19635 ( .A0(n9834), .A1(n9828), .S(n4131), .Z(n9841) );
  CMX2X1 U19636 ( .A0(n9829), .A1(n9841), .S(n3797), .Z(n9854) );
  CMXI2X1 U19637 ( .A0(n9830), .A1(n9854), .S(n3505), .Z(N5309) );
  CMX2X1 U19638 ( .A0(N8113), .A1(N8112), .S(n4280), .Z(n9837) );
  CMXI2X1 U19639 ( .A0(n9837), .A1(n9831), .S(n4131), .Z(n9844) );
  CMX2X1 U19640 ( .A0(n9832), .A1(n9844), .S(n3805), .Z(n9861) );
  CMXI2X1 U19641 ( .A0(n9833), .A1(n9861), .S(n3505), .Z(N5310) );
  CMX2X1 U19642 ( .A0(N8112), .A1(N8111), .S(n4280), .Z(n9840) );
  CMXI2X1 U19643 ( .A0(n9840), .A1(n9834), .S(n4131), .Z(n9847) );
  CMX2X1 U19644 ( .A0(n9835), .A1(n9847), .S(n3806), .Z(n9864) );
  CMXI2X1 U19645 ( .A0(n9836), .A1(n9864), .S(n3505), .Z(N5311) );
  CMX2X1 U19646 ( .A0(N8111), .A1(N8110), .S(n4280), .Z(n9843) );
  CMXI2X1 U19647 ( .A0(n9843), .A1(n9837), .S(n4131), .Z(n9850) );
  CMX2X1 U19648 ( .A0(n9838), .A1(n9850), .S(n3807), .Z(n9867) );
  CMXI2X1 U19649 ( .A0(n9839), .A1(n9867), .S(n3504), .Z(N5312) );
  CMX2X1 U19650 ( .A0(N8110), .A1(N8109), .S(n4279), .Z(n9846) );
  CMXI2X1 U19651 ( .A0(n9846), .A1(n9840), .S(n4131), .Z(n9853) );
  CMX2X1 U19652 ( .A0(n9841), .A1(n9853), .S(n3808), .Z(n9870) );
  CMXI2X1 U19653 ( .A0(n9842), .A1(n9870), .S(n3504), .Z(N5313) );
  CMX2X1 U19654 ( .A0(N8109), .A1(N8108), .S(n4279), .Z(n9849) );
  CMXI2X1 U19655 ( .A0(n9849), .A1(n9843), .S(n4131), .Z(n9860) );
  CMX2X1 U19656 ( .A0(n9844), .A1(n9860), .S(n3808), .Z(n9873) );
  CMXI2X1 U19657 ( .A0(n9845), .A1(n9873), .S(n3504), .Z(N5314) );
  CMX2X1 U19658 ( .A0(N8108), .A1(N8107), .S(n4279), .Z(n9852) );
  CMXI2X1 U19659 ( .A0(n9852), .A1(n9846), .S(n4131), .Z(n9863) );
  CMX2X1 U19660 ( .A0(n9847), .A1(n9863), .S(n3772), .Z(n9876) );
  CMXI2X1 U19661 ( .A0(n9848), .A1(n9876), .S(n3508), .Z(N5315) );
  CMX2X1 U19662 ( .A0(N8107), .A1(N8106), .S(n4279), .Z(n9859) );
  CMXI2X1 U19663 ( .A0(n9859), .A1(n9849), .S(n4131), .Z(n9866) );
  CMX2X1 U19664 ( .A0(n9850), .A1(n9866), .S(n3773), .Z(n9879) );
  CMXI2X1 U19665 ( .A0(n9851), .A1(n9879), .S(n3507), .Z(N5316) );
  CMX2X1 U19666 ( .A0(N8106), .A1(N8105), .S(n4279), .Z(n9862) );
  CMXI2X1 U19667 ( .A0(n9862), .A1(n9852), .S(n4131), .Z(n9869) );
  CMX2X1 U19668 ( .A0(n9853), .A1(n9869), .S(n3774), .Z(n9882) );
  CMXI2X1 U19669 ( .A0(n9854), .A1(n9882), .S(n3507), .Z(N5317) );
  CMX2X1 U19670 ( .A0(n9856), .A1(n9855), .S(n3775), .Z(n12006) );
  CMX2X1 U19671 ( .A0(N8250), .A1(N8249), .S(n4279), .Z(n9925) );
  CMXI2X1 U19672 ( .A0(n9925), .A1(n9857), .S(n4131), .Z(n9991) );
  CMX2X1 U19673 ( .A0(n9858), .A1(n9991), .S(n3776), .Z(n10129) );
  CMXI2X1 U19674 ( .A0(n12006), .A1(n10129), .S(n3507), .Z(N5173) );
  CMX2X1 U19675 ( .A0(N8105), .A1(N8104), .S(n4279), .Z(n9865) );
  CMXI2X1 U19676 ( .A0(n9865), .A1(n9859), .S(n4131), .Z(n9872) );
  CMX2X1 U19677 ( .A0(n9860), .A1(n9872), .S(n3777), .Z(n9885) );
  CMXI2X1 U19678 ( .A0(n9861), .A1(n9885), .S(n3507), .Z(N5318) );
  CMX2X1 U19679 ( .A0(N8104), .A1(N8103), .S(n4279), .Z(n9868) );
  CMXI2X1 U19680 ( .A0(n9868), .A1(n9862), .S(n4130), .Z(n9875) );
  CMX2X1 U19681 ( .A0(n9863), .A1(n9875), .S(n3790), .Z(n9888) );
  CMXI2X1 U19682 ( .A0(n9864), .A1(n9888), .S(n3507), .Z(N5319) );
  CMX2X1 U19683 ( .A0(N8103), .A1(N8102), .S(n4279), .Z(n9871) );
  CMXI2X1 U19684 ( .A0(n9871), .A1(n9865), .S(n4130), .Z(n9878) );
  CMX2X1 U19685 ( .A0(n9866), .A1(n9878), .S(n3793), .Z(n9895) );
  CMXI2X1 U19686 ( .A0(n9867), .A1(n9895), .S(n3507), .Z(N5320) );
  CMX2X1 U19687 ( .A0(N8102), .A1(N8101), .S(n4279), .Z(n9874) );
  CMXI2X1 U19688 ( .A0(n9874), .A1(n9868), .S(n4130), .Z(n9881) );
  CMX2X1 U19689 ( .A0(n9869), .A1(n9881), .S(n3794), .Z(n9898) );
  CMXI2X1 U19690 ( .A0(n9870), .A1(n9898), .S(n3507), .Z(N5321) );
  CMX2X1 U19691 ( .A0(N8101), .A1(N8100), .S(n4279), .Z(n9877) );
  CMXI2X1 U19692 ( .A0(n9877), .A1(n9871), .S(n4130), .Z(n9884) );
  CMX2X1 U19693 ( .A0(n9872), .A1(n9884), .S(n3795), .Z(n9901) );
  CMXI2X1 U19694 ( .A0(n9873), .A1(n9901), .S(n3507), .Z(N5322) );
  CMX2X1 U19695 ( .A0(N8100), .A1(N8099), .S(n4278), .Z(n9880) );
  CMXI2X1 U19696 ( .A0(n9880), .A1(n9874), .S(n4130), .Z(n9887) );
  CMX2X1 U19697 ( .A0(n9875), .A1(n9887), .S(n3796), .Z(n9904) );
  CMXI2X1 U19698 ( .A0(n9876), .A1(n9904), .S(n3507), .Z(N5323) );
  CMX2X1 U19699 ( .A0(N8099), .A1(N8098), .S(n4278), .Z(n9883) );
  CMXI2X1 U19700 ( .A0(n9883), .A1(n9877), .S(n4130), .Z(n9894) );
  CMX2X1 U19701 ( .A0(n9878), .A1(n9894), .S(n3797), .Z(n9907) );
  CMXI2X1 U19702 ( .A0(n9879), .A1(n9907), .S(n3507), .Z(N5324) );
  CMX2X1 U19703 ( .A0(N8098), .A1(N8097), .S(n4278), .Z(n9886) );
  CMXI2X1 U19704 ( .A0(n9886), .A1(n9880), .S(n4130), .Z(n9897) );
  CMX2X1 U19705 ( .A0(n9881), .A1(n9897), .S(n3805), .Z(n9910) );
  CMXI2X1 U19706 ( .A0(n9882), .A1(n9910), .S(n3506), .Z(N5325) );
  CMX2X1 U19707 ( .A0(N8097), .A1(N8096), .S(n4281), .Z(n9893) );
  CMXI2X1 U19708 ( .A0(n9893), .A1(n9883), .S(n4130), .Z(n9900) );
  CMX2X1 U19709 ( .A0(n9884), .A1(n9900), .S(n3806), .Z(n9913) );
  CMXI2X1 U19710 ( .A0(n9885), .A1(n9913), .S(n3506), .Z(N5326) );
  CMX2X1 U19711 ( .A0(N8096), .A1(N8095), .S(n4250), .Z(n9896) );
  CMXI2X1 U19712 ( .A0(n9896), .A1(n9886), .S(n4130), .Z(n9903) );
  CMX2X1 U19713 ( .A0(n9887), .A1(n9903), .S(n3807), .Z(n9916) );
  CMXI2X1 U19714 ( .A0(n9888), .A1(n9916), .S(n3506), .Z(N5327) );
  CMX2X1 U19715 ( .A0(n9890), .A1(n9889), .S(n3808), .Z(n12340) );
  CMX2X1 U19716 ( .A0(N8249), .A1(N8248), .S(n4250), .Z(n9957) );
  CMXI2X1 U19717 ( .A0(n9957), .A1(n9891), .S(n4130), .Z(n10029) );
  CMX2X1 U19718 ( .A0(n9892), .A1(n10029), .S(n3809), .Z(n10162) );
  CMXI2X1 U19719 ( .A0(n12340), .A1(n10162), .S(n3506), .Z(N5174) );
  CMX2X1 U19720 ( .A0(N8095), .A1(N8094), .S(n4249), .Z(n9899) );
  CMXI2X1 U19721 ( .A0(n9899), .A1(n9893), .S(n4130), .Z(n9906) );
  CMX2X1 U19722 ( .A0(n9894), .A1(n9906), .S(n3810), .Z(n9919) );
  CMXI2X1 U19723 ( .A0(n9895), .A1(n9919), .S(n3506), .Z(N5328) );
  CMX2X1 U19724 ( .A0(N8094), .A1(N8093), .S(n4249), .Z(n9902) );
  CMXI2X1 U19725 ( .A0(n9902), .A1(n9896), .S(n4130), .Z(n9909) );
  CMX2X1 U19726 ( .A0(n9897), .A1(n9909), .S(n3811), .Z(n9922) );
  CMXI2X1 U19727 ( .A0(n9898), .A1(n9922), .S(n3506), .Z(N5329) );
  CMX2X1 U19728 ( .A0(N8093), .A1(N8092), .S(n4249), .Z(n9905) );
  CMXI2X1 U19729 ( .A0(n9905), .A1(n9899), .S(n4130), .Z(n9912) );
  CMX2X1 U19730 ( .A0(n9900), .A1(n9912), .S(n3812), .Z(n9929) );
  CMXI2X1 U19731 ( .A0(n9901), .A1(n9929), .S(n3506), .Z(N5330) );
  CMX2X1 U19732 ( .A0(N8092), .A1(N8091), .S(n4249), .Z(n9908) );
  CMXI2X1 U19733 ( .A0(n9908), .A1(n9902), .S(n4130), .Z(n9915) );
  CMX2X1 U19734 ( .A0(n9903), .A1(n9915), .S(n4326), .Z(n9932) );
  CMXI2X1 U19735 ( .A0(n9904), .A1(n9932), .S(n3509), .Z(N5331) );
  CMXI2X1 U19736 ( .A0(n9911), .A1(n9905), .S(n4130), .Z(n9918) );
  CMX2X1 U19737 ( .A0(n9906), .A1(n9918), .S(n3771), .Z(n9935) );
  CMXI2X1 U19738 ( .A0(n9907), .A1(n9935), .S(n3509), .Z(N5332) );
  CMXI2X1 U19739 ( .A0(n9914), .A1(n9908), .S(n4130), .Z(n9921) );
  CMX2X1 U19740 ( .A0(n9909), .A1(n9921), .S(n3808), .Z(n9938) );
  CMXI2X1 U19741 ( .A0(n9910), .A1(n9938), .S(n3509), .Z(N5333) );
  CMX2X1 U19742 ( .A0(N8089), .A1(N8088), .S(n4249), .Z(n9917) );
  CMXI2X1 U19743 ( .A0(n9917), .A1(n9911), .S(n4129), .Z(n9928) );
  CMX2X1 U19744 ( .A0(n9912), .A1(n9928), .S(n3809), .Z(n9941) );
  CMXI2X1 U19745 ( .A0(n9913), .A1(n9941), .S(n3509), .Z(N5334) );
  CMX2X1 U19746 ( .A0(N8088), .A1(N8087), .S(n4249), .Z(n9920) );
  CMXI2X1 U19747 ( .A0(n9920), .A1(n9914), .S(n4129), .Z(n9931) );
  CMX2X1 U19748 ( .A0(n9915), .A1(n9931), .S(n3792), .Z(n9944) );
  CMXI2X1 U19749 ( .A0(n9916), .A1(n9944), .S(n3509), .Z(N5335) );
  CMX2X1 U19750 ( .A0(N8087), .A1(N8086), .S(n4249), .Z(n9927) );
  CMXI2X1 U19751 ( .A0(n9927), .A1(n9917), .S(n4129), .Z(n9934) );
  CMX2X1 U19752 ( .A0(n9918), .A1(n9934), .S(n3793), .Z(n9947) );
  CMXI2X1 U19753 ( .A0(n9919), .A1(n9947), .S(n3509), .Z(N5336) );
  CMX2X1 U19754 ( .A0(N8086), .A1(N8085), .S(n4249), .Z(n9930) );
  CMXI2X1 U19755 ( .A0(n9930), .A1(n9920), .S(n4129), .Z(n9937) );
  CMX2X1 U19756 ( .A0(n9921), .A1(n9937), .S(n3794), .Z(n9950) );
  CMXI2X1 U19757 ( .A0(n9922), .A1(n9950), .S(n3509), .Z(N5337) );
  CMX2X1 U19758 ( .A0(n9924), .A1(n9923), .S(n3795), .Z(n12658) );
  CMX2X1 U19759 ( .A0(N8248), .A1(N8247), .S(n4249), .Z(n9990) );
  CMXI2X1 U19760 ( .A0(n9990), .A1(n9925), .S(n4129), .Z(n10062) );
  CMX2X1 U19761 ( .A0(n9926), .A1(n10062), .S(n3796), .Z(n10195) );
  CMXI2X1 U19762 ( .A0(n12658), .A1(n10195), .S(n3509), .Z(N5175) );
  CMX2X1 U19763 ( .A0(N8085), .A1(N8084), .S(n4248), .Z(n9933) );
  CMXI2X1 U19764 ( .A0(n9933), .A1(n9927), .S(n4129), .Z(n9940) );
  CMX2X1 U19765 ( .A0(n9928), .A1(n9940), .S(n3805), .Z(n9953) );
  CMXI2X1 U19766 ( .A0(n9929), .A1(n9953), .S(n3508), .Z(N5338) );
  CMX2X1 U19767 ( .A0(N8084), .A1(N8083), .S(n4248), .Z(n9936) );
  CMXI2X1 U19768 ( .A0(n9936), .A1(n9930), .S(n4129), .Z(n9943) );
  CMX2X1 U19769 ( .A0(n9931), .A1(n9943), .S(n3806), .Z(n9956) );
  CMXI2X1 U19770 ( .A0(n9932), .A1(n9956), .S(n3508), .Z(N5339) );
  CMX2X1 U19771 ( .A0(N8083), .A1(N8082), .S(n4248), .Z(n9939) );
  CMXI2X1 U19772 ( .A0(n9939), .A1(n9933), .S(n4129), .Z(n9946) );
  CMX2X1 U19773 ( .A0(n9934), .A1(n9946), .S(n3808), .Z(n9962) );
  CMXI2X1 U19774 ( .A0(n9935), .A1(n9962), .S(n3508), .Z(N5340) );
  CMX2X1 U19775 ( .A0(N8082), .A1(N8081), .S(n4248), .Z(n9942) );
  CMXI2X1 U19776 ( .A0(n9942), .A1(n9936), .S(n4129), .Z(n9949) );
  CMX2X1 U19777 ( .A0(n9937), .A1(n9949), .S(n3809), .Z(n9965) );
  CMXI2X1 U19778 ( .A0(n9938), .A1(n9965), .S(n3508), .Z(N5341) );
  CMX2X1 U19779 ( .A0(N8081), .A1(N8080), .S(n4248), .Z(n9945) );
  CMXI2X1 U19780 ( .A0(n9945), .A1(n9939), .S(n4129), .Z(n9952) );
  CMX2X1 U19781 ( .A0(n9940), .A1(n9952), .S(n3810), .Z(n9968) );
  CMXI2X1 U19782 ( .A0(n9941), .A1(n9968), .S(n3508), .Z(N5342) );
  CMX2X1 U19783 ( .A0(N8080), .A1(N8079), .S(n4248), .Z(n9948) );
  CMXI2X1 U19784 ( .A0(n9948), .A1(n9942), .S(n4129), .Z(n9955) );
  CMX2X1 U19785 ( .A0(n9943), .A1(n9955), .S(n3797), .Z(n9971) );
  CMXI2X1 U19786 ( .A0(n9944), .A1(n9971), .S(n3508), .Z(N5343) );
  CMX2X1 U19787 ( .A0(N8079), .A1(N8078), .S(n4248), .Z(n9951) );
  CMXI2X1 U19788 ( .A0(n9951), .A1(n9945), .S(n4129), .Z(n9961) );
  CMX2X1 U19789 ( .A0(n9946), .A1(n9961), .S(n3805), .Z(n9974) );
  CMXI2X1 U19790 ( .A0(n9947), .A1(n9974), .S(n3508), .Z(N5344) );
  CMX2X1 U19791 ( .A0(N8078), .A1(N8077), .S(n4248), .Z(n9954) );
  CMXI2X1 U19792 ( .A0(n9954), .A1(n9948), .S(n4129), .Z(n9964) );
  CMX2X1 U19793 ( .A0(n9949), .A1(n9964), .S(n3806), .Z(n9977) );
  CMXI2X1 U19794 ( .A0(n9950), .A1(n9977), .S(n3508), .Z(N5345) );
  CMX2X1 U19795 ( .A0(N8077), .A1(N8076), .S(n4248), .Z(n9960) );
  CMXI2X1 U19796 ( .A0(n9960), .A1(n9951), .S(n4129), .Z(n9967) );
  CMX2X1 U19797 ( .A0(n9952), .A1(n9967), .S(n4307), .Z(n9980) );
  CMXI2X1 U19798 ( .A0(n9953), .A1(n9980), .S(n3508), .Z(N5346) );
  CMX2X1 U19799 ( .A0(N8076), .A1(N8075), .S(n4248), .Z(n9963) );
  CMXI2X1 U19800 ( .A0(n9963), .A1(n9954), .S(n4129), .Z(n9970) );
  CMX2X1 U19801 ( .A0(n9955), .A1(n9970), .S(n3806), .Z(n9983) );
  CMXI2X1 U19802 ( .A0(n9956), .A1(n9983), .S(n3508), .Z(N5347) );
  CMX2X1 U19803 ( .A0(N8247), .A1(N8246), .S(n4248), .Z(n10028) );
  CMXI2X1 U19804 ( .A0(n10028), .A1(n9957), .S(n4129), .Z(n10095) );
  CMX2X1 U19805 ( .A0(n9958), .A1(n10095), .S(n3775), .Z(n10228) );
  CMXI2X1 U19806 ( .A0(n9959), .A1(n10228), .S(n3317), .Z(N5176) );
  CMX2X1 U19807 ( .A0(N8075), .A1(N8074), .S(n4247), .Z(n9966) );
  CMXI2X1 U19808 ( .A0(n9966), .A1(n9960), .S(n4128), .Z(n9973) );
  CMX2X1 U19809 ( .A0(n9961), .A1(n9973), .S(n3776), .Z(n9986) );
  CMXI2X1 U19810 ( .A0(n9962), .A1(n9986), .S(n3317), .Z(N5348) );
  CMX2X1 U19811 ( .A0(N8074), .A1(N8073), .S(n4247), .Z(n9969) );
  CMXI2X1 U19812 ( .A0(n9969), .A1(n9963), .S(n4128), .Z(n9976) );
  CMX2X1 U19813 ( .A0(n9964), .A1(n9976), .S(n3777), .Z(n9989) );
  CMXI2X1 U19814 ( .A0(n9965), .A1(n9989), .S(n3317), .Z(N5349) );
  CMX2X1 U19815 ( .A0(N8073), .A1(N8072), .S(n4247), .Z(n9972) );
  CMXI2X1 U19816 ( .A0(n9972), .A1(n9966), .S(n4128), .Z(n9979) );
  CMX2X1 U19817 ( .A0(n9967), .A1(n9979), .S(n3790), .Z(n10000) );
  CMXI2X1 U19818 ( .A0(n9968), .A1(n10000), .S(n3396), .Z(N5350) );
  CMX2X1 U19819 ( .A0(N8072), .A1(N8071), .S(n4247), .Z(n9975) );
  CMXI2X1 U19820 ( .A0(n9975), .A1(n9969), .S(n4128), .Z(n9982) );
  CMX2X1 U19821 ( .A0(n9970), .A1(n9982), .S(n3791), .Z(n10003) );
  CMXI2X1 U19822 ( .A0(n9971), .A1(n10003), .S(n3423), .Z(N5351) );
  CMX2X1 U19823 ( .A0(N8071), .A1(N8070), .S(n4247), .Z(n9978) );
  CMXI2X1 U19824 ( .A0(n9978), .A1(n9972), .S(n4128), .Z(n9985) );
  CMX2X1 U19825 ( .A0(n9973), .A1(n9985), .S(n3806), .Z(n10006) );
  CMXI2X1 U19826 ( .A0(n9974), .A1(n10006), .S(n3423), .Z(N5352) );
  CMX2X1 U19827 ( .A0(N8070), .A1(N8069), .S(n4247), .Z(n9981) );
  CMXI2X1 U19828 ( .A0(n9981), .A1(n9975), .S(n4128), .Z(n9988) );
  CMX2X1 U19829 ( .A0(n9976), .A1(n9988), .S(n3807), .Z(n10009) );
  CMXI2X1 U19830 ( .A0(n9977), .A1(n10009), .S(n3423), .Z(N5353) );
  CMX2X1 U19831 ( .A0(N8069), .A1(N8068), .S(n4247), .Z(n9984) );
  CMXI2X1 U19832 ( .A0(n9984), .A1(n9978), .S(n4128), .Z(n9999) );
  CMX2X1 U19833 ( .A0(n9979), .A1(n9999), .S(n3808), .Z(n10012) );
  CMXI2X1 U19834 ( .A0(n9980), .A1(n10012), .S(n3423), .Z(N5354) );
  CMX2X1 U19835 ( .A0(N8068), .A1(N8067), .S(n4247), .Z(n9987) );
  CMXI2X1 U19836 ( .A0(n9987), .A1(n9981), .S(n4128), .Z(n10002) );
  CMX2X1 U19837 ( .A0(n9982), .A1(n10002), .S(n3809), .Z(n10015) );
  CMXI2X1 U19838 ( .A0(n9983), .A1(n10015), .S(n3423), .Z(N5355) );
  CMX2X1 U19839 ( .A0(N8067), .A1(N8066), .S(n4247), .Z(n9998) );
  CMXI2X1 U19840 ( .A0(n9998), .A1(n9984), .S(n4128), .Z(n10005) );
  CMX2X1 U19841 ( .A0(n9985), .A1(n10005), .S(n3810), .Z(n10018) );
  CMXI2X1 U19842 ( .A0(n9986), .A1(n10018), .S(n3423), .Z(N5356) );
  CMX2X1 U19843 ( .A0(N8066), .A1(N8065), .S(n4247), .Z(n10001) );
  CMXI2X1 U19844 ( .A0(n10001), .A1(n9987), .S(n4128), .Z(n10008) );
  CMX2X1 U19845 ( .A0(n9988), .A1(n10008), .S(n3811), .Z(n10021) );
  CMXI2X1 U19846 ( .A0(n9989), .A1(n10021), .S(n3422), .Z(N5357) );
  CMX2X1 U19847 ( .A0(N8246), .A1(N8245), .S(n4247), .Z(n10061) );
  CMXI2X1 U19848 ( .A0(n10061), .A1(n9990), .S(n4128), .Z(n10128) );
  CMX2X1 U19849 ( .A0(n9991), .A1(n10128), .S(n3812), .Z(n10261) );
  CMXI2X1 U19850 ( .A0(n9992), .A1(n10261), .S(n3422), .Z(N5177) );
  CMXI2X1 U19851 ( .A0(N8271), .A1(N8272), .S(n3883), .Z(n10665) );
  CMXI2X1 U19852 ( .A0(N8273), .A1(N8274), .S(n3885), .Z(n10668) );
  CMXI2X1 U19853 ( .A0(n10665), .A1(n10668), .S(n4128), .Z(n11337) );
  CMXI2X1 U19854 ( .A0(N8276), .A1(N8275), .S(n3868), .Z(n10667) );
  CMXI2X1 U19855 ( .A0(N8277), .A1(N8278), .S(n3887), .Z(n9993) );
  CMXI2X1 U19856 ( .A0(n10667), .A1(n9993), .S(n4128), .Z(n9994) );
  CMXI2X1 U19857 ( .A0(n11337), .A1(n9994), .S(n3783), .Z(n9997) );
  CMXI2X1 U19858 ( .A0(N8269), .A1(N8270), .S(n3887), .Z(n10666) );
  CMXI2X1 U19859 ( .A0(n9995), .A1(n4431), .S(n4128), .Z(n11336) );
  CMX2X1 U19860 ( .A0(n11336), .A1(n9996), .S(n4312), .Z(n12659) );
  CMXI2X1 U19861 ( .A0(n9997), .A1(n12659), .S(n3422), .Z(N5159) );
  CMX2X1 U19862 ( .A0(N8065), .A1(N8064), .S(n4246), .Z(n10004) );
  CMXI2X1 U19863 ( .A0(n10004), .A1(n9998), .S(n4128), .Z(n10011) );
  CMX2X1 U19864 ( .A0(n9999), .A1(n10011), .S(n3771), .Z(n10024) );
  CMXI2X1 U19865 ( .A0(n10000), .A1(n10024), .S(n3422), .Z(N5358) );
  CMX2X1 U19866 ( .A0(N8064), .A1(N8063), .S(n4246), .Z(n10007) );
  CMXI2X1 U19867 ( .A0(n10007), .A1(n10001), .S(n4128), .Z(n10014) );
  CMX2X1 U19868 ( .A0(n10002), .A1(n10014), .S(n3772), .Z(n10027) );
  CMXI2X1 U19869 ( .A0(n10003), .A1(n10027), .S(n3422), .Z(N5359) );
  CMX2X1 U19870 ( .A0(N8063), .A1(N8062), .S(n4246), .Z(n10010) );
  CMXI2X1 U19871 ( .A0(n10010), .A1(n10004), .S(n4127), .Z(n10017) );
  CMX2X1 U19872 ( .A0(n10005), .A1(n10017), .S(n3773), .Z(n10033) );
  CMXI2X1 U19873 ( .A0(n10006), .A1(n10033), .S(n3422), .Z(N5360) );
  CMX2X1 U19874 ( .A0(N8062), .A1(N8061), .S(n4246), .Z(n10013) );
  CMXI2X1 U19875 ( .A0(n10013), .A1(n10007), .S(n4127), .Z(n10020) );
  CMX2X1 U19876 ( .A0(n10008), .A1(n10020), .S(n3774), .Z(n10036) );
  CMXI2X1 U19877 ( .A0(n10009), .A1(n10036), .S(n3422), .Z(N5361) );
  CMX2X1 U19878 ( .A0(N8061), .A1(N8060), .S(n4246), .Z(n10016) );
  CMXI2X1 U19879 ( .A0(n10016), .A1(n10010), .S(n4127), .Z(n10023) );
  CMX2X1 U19880 ( .A0(n10011), .A1(n10023), .S(n3807), .Z(n10039) );
  CMXI2X1 U19881 ( .A0(n10012), .A1(n10039), .S(n3422), .Z(N5362) );
  CMX2X1 U19882 ( .A0(N8060), .A1(N8059), .S(n4246), .Z(n10019) );
  CMXI2X1 U19883 ( .A0(n10019), .A1(n10013), .S(n4127), .Z(n10026) );
  CMX2X1 U19884 ( .A0(n10014), .A1(n10026), .S(n3808), .Z(n10042) );
  CMXI2X1 U19885 ( .A0(n10015), .A1(n10042), .S(n3422), .Z(N5363) );
  CMX2X1 U19886 ( .A0(N8059), .A1(N8058), .S(n4246), .Z(n10022) );
  CMXI2X1 U19887 ( .A0(n10022), .A1(n10016), .S(n4127), .Z(n10032) );
  CMX2X1 U19888 ( .A0(n10017), .A1(n10032), .S(n3809), .Z(n10045) );
  CMXI2X1 U19889 ( .A0(n10018), .A1(n10045), .S(n3425), .Z(N5364) );
  CMXI2X1 U19890 ( .A0(n10025), .A1(n10019), .S(n4127), .Z(n10035) );
  CMX2X1 U19891 ( .A0(n10020), .A1(n10035), .S(n3810), .Z(n10048) );
  CMXI2X1 U19892 ( .A0(n10021), .A1(n10048), .S(n3425), .Z(N5365) );
  CMX2X1 U19893 ( .A0(N8057), .A1(N8056), .S(n4246), .Z(n10031) );
  CMXI2X1 U19894 ( .A0(n10031), .A1(n10022), .S(n4127), .Z(n10038) );
  CMX2X1 U19895 ( .A0(n10023), .A1(n10038), .S(n3809), .Z(n10051) );
  CMXI2X1 U19896 ( .A0(n10024), .A1(n10051), .S(n3425), .Z(N5366) );
  CMX2X1 U19897 ( .A0(N8056), .A1(N8055), .S(n4246), .Z(n10034) );
  CMXI2X1 U19898 ( .A0(n10034), .A1(n10025), .S(n4127), .Z(n10041) );
  CMX2X1 U19899 ( .A0(n10026), .A1(n10041), .S(n3792), .Z(n10054) );
  CMXI2X1 U19900 ( .A0(n10027), .A1(n10054), .S(n3425), .Z(N5367) );
  CMXI2X1 U19901 ( .A0(n10094), .A1(n10028), .S(n4127), .Z(n10161) );
  CMX2X1 U19902 ( .A0(n10029), .A1(n10161), .S(n3793), .Z(n10294) );
  CMXI2X1 U19903 ( .A0(n10030), .A1(n10294), .S(n3425), .Z(N5178) );
  CMX2X1 U19904 ( .A0(N8055), .A1(N8054), .S(n4245), .Z(n10037) );
  CMXI2X1 U19905 ( .A0(n10037), .A1(n10031), .S(n4127), .Z(n10044) );
  CMX2X1 U19906 ( .A0(n10032), .A1(n10044), .S(n3794), .Z(n10057) );
  CMXI2X1 U19907 ( .A0(n10033), .A1(n10057), .S(n3424), .Z(N5368) );
  CMX2X1 U19908 ( .A0(N8054), .A1(N8053), .S(n4245), .Z(n10040) );
  CMXI2X1 U19909 ( .A0(n10040), .A1(n10034), .S(n4127), .Z(n10047) );
  CMX2X1 U19910 ( .A0(n10035), .A1(n10047), .S(n3795), .Z(n10060) );
  CMXI2X1 U19911 ( .A0(n10036), .A1(n10060), .S(n3424), .Z(N5369) );
  CMXI2X1 U19912 ( .A0(n10043), .A1(n10037), .S(n4127), .Z(n10050) );
  CMX2X1 U19913 ( .A0(n10038), .A1(n10050), .S(n3796), .Z(n10066) );
  CMXI2X1 U19914 ( .A0(n10039), .A1(n10066), .S(n3424), .Z(N5370) );
  CMXI2X1 U19915 ( .A0(n10046), .A1(n10040), .S(n4127), .Z(n10053) );
  CMX2X1 U19916 ( .A0(n10041), .A1(n10053), .S(n3797), .Z(n10069) );
  CMXI2X1 U19917 ( .A0(n10042), .A1(n10069), .S(n3424), .Z(N5371) );
  CMXI2X1 U19918 ( .A0(n10049), .A1(n10043), .S(n4127), .Z(n10056) );
  CMX2X1 U19919 ( .A0(n10044), .A1(n10056), .S(n3805), .Z(n10072) );
  CMXI2X1 U19920 ( .A0(n10045), .A1(n10072), .S(n3424), .Z(N5372) );
  CMXI2X1 U19921 ( .A0(n10052), .A1(n10046), .S(n4127), .Z(n10059) );
  CMX2X1 U19922 ( .A0(n10047), .A1(n10059), .S(n3806), .Z(n10075) );
  CMXI2X1 U19923 ( .A0(n10048), .A1(n10075), .S(n3424), .Z(N5373) );
  CMXI2X1 U19924 ( .A0(n10055), .A1(n10049), .S(n4127), .Z(n10065) );
  CMX2X1 U19925 ( .A0(n10050), .A1(n10065), .S(n3807), .Z(n10078) );
  CMXI2X1 U19926 ( .A0(n10051), .A1(n10078), .S(n3424), .Z(N5374) );
  CMXI2X1 U19927 ( .A0(n10058), .A1(n10052), .S(n4126), .Z(n10068) );
  CMX2X1 U19928 ( .A0(n10053), .A1(n10068), .S(n3808), .Z(n10081) );
  CMXI2X1 U19929 ( .A0(n10054), .A1(n10081), .S(n3424), .Z(N5375) );
  CMXI2X1 U19930 ( .A0(n10064), .A1(n10055), .S(n4126), .Z(n10071) );
  CMX2X1 U19931 ( .A0(n10056), .A1(n10071), .S(n3809), .Z(n10084) );
  CMXI2X1 U19932 ( .A0(n10057), .A1(n10084), .S(n3424), .Z(N5376) );
  CMX2X1 U19933 ( .A0(N8046), .A1(N8045), .S(n4245), .Z(n10067) );
  CMXI2X1 U19934 ( .A0(n10067), .A1(n10058), .S(n4126), .Z(n10074) );
  CMX2X1 U19935 ( .A0(n10059), .A1(n10074), .S(n3810), .Z(n10087) );
  CMXI2X1 U19936 ( .A0(n10060), .A1(n10087), .S(n3424), .Z(N5377) );
  CMXI2X1 U19937 ( .A0(n10127), .A1(n10061), .S(n4126), .Z(n10194) );
  CMX2X1 U19938 ( .A0(n10062), .A1(n10194), .S(n3811), .Z(n10327) );
  CMXI2X1 U19939 ( .A0(n10063), .A1(n10327), .S(n3424), .Z(N5179) );
  CMX2X1 U19940 ( .A0(N8045), .A1(N8044), .S(n4244), .Z(n10070) );
  CMXI2X1 U19941 ( .A0(n10070), .A1(n10064), .S(n4126), .Z(n10077) );
  CMX2X1 U19942 ( .A0(n10065), .A1(n10077), .S(n3812), .Z(n10090) );
  CMXI2X1 U19943 ( .A0(n10066), .A1(n10090), .S(n3423), .Z(N5378) );
  CMX2X1 U19944 ( .A0(N8044), .A1(N8043), .S(n4244), .Z(n10073) );
  CMXI2X1 U19945 ( .A0(n10073), .A1(n10067), .S(n4126), .Z(n10080) );
  CMX2X1 U19946 ( .A0(n10068), .A1(n10080), .S(n4336), .Z(n10093) );
  CMXI2X1 U19947 ( .A0(n10069), .A1(n10093), .S(n3423), .Z(N5379) );
  CMX2X1 U19948 ( .A0(N8043), .A1(N8042), .S(n4244), .Z(n10076) );
  CMXI2X1 U19949 ( .A0(n10076), .A1(n10070), .S(n4126), .Z(n10083) );
  CMX2X1 U19950 ( .A0(n10071), .A1(n10083), .S(n3771), .Z(n10099) );
  CMXI2X1 U19951 ( .A0(n10072), .A1(n10099), .S(n3427), .Z(N5380) );
  CMXI2X1 U19952 ( .A0(n10079), .A1(n10073), .S(n4126), .Z(n10086) );
  CMX2X1 U19953 ( .A0(n10074), .A1(n10086), .S(n3777), .Z(n10102) );
  CMXI2X1 U19954 ( .A0(n10075), .A1(n10102), .S(n3426), .Z(N5381) );
  CMXI2X1 U19955 ( .A0(n10082), .A1(n10076), .S(n4126), .Z(n10089) );
  CMX2X1 U19956 ( .A0(n10077), .A1(n10089), .S(n3790), .Z(n10105) );
  CMXI2X1 U19957 ( .A0(n10078), .A1(n10105), .S(n3426), .Z(N5382) );
  CMXI2X1 U19958 ( .A0(n10085), .A1(n10079), .S(n4126), .Z(n10092) );
  CMX2X1 U19959 ( .A0(n10080), .A1(n10092), .S(n3811), .Z(n10108) );
  CMXI2X1 U19960 ( .A0(n10081), .A1(n10108), .S(n3426), .Z(N5383) );
  CMXI2X1 U19961 ( .A0(n10088), .A1(n10082), .S(n4126), .Z(n10098) );
  CMX2X1 U19962 ( .A0(n10083), .A1(n10098), .S(n3812), .Z(n10111) );
  CMXI2X1 U19963 ( .A0(n10084), .A1(n10111), .S(n3426), .Z(N5384) );
  CMXI2X1 U19964 ( .A0(n10091), .A1(n10085), .S(n4126), .Z(n10101) );
  CMX2X1 U19965 ( .A0(n10086), .A1(n10101), .S(n4307), .Z(n10114) );
  CMXI2X1 U19966 ( .A0(n10087), .A1(n10114), .S(n3426), .Z(N5385) );
  CMXI2X1 U19967 ( .A0(n10097), .A1(n10088), .S(n4126), .Z(n10104) );
  CMX2X1 U19968 ( .A0(n10089), .A1(n10104), .S(n3771), .Z(n10117) );
  CMXI2X1 U19969 ( .A0(n10090), .A1(n10117), .S(n3426), .Z(N5386) );
  CMXI2X1 U19970 ( .A0(n10100), .A1(n10091), .S(n4126), .Z(n10107) );
  CMX2X1 U19971 ( .A0(n10092), .A1(n10107), .S(n3772), .Z(n10120) );
  CMXI2X1 U19972 ( .A0(n10093), .A1(n10120), .S(n3426), .Z(N5387) );
  CMX2X1 U19973 ( .A0(N8243), .A1(N8242), .S(n4244), .Z(n10160) );
  CMXI2X1 U19974 ( .A0(n10160), .A1(n10094), .S(n4126), .Z(n10227) );
  CMX2X1 U19975 ( .A0(n10095), .A1(n10227), .S(n3810), .Z(n10367) );
  CMXI2X1 U19976 ( .A0(n10096), .A1(n10367), .S(n3426), .Z(N5180) );
  CMXI2X1 U19977 ( .A0(n10103), .A1(n10097), .S(n4126), .Z(n10110) );
  CMX2X1 U19978 ( .A0(n10098), .A1(n10110), .S(n3772), .Z(n10123) );
  CMXI2X1 U19979 ( .A0(n10099), .A1(n10123), .S(n3426), .Z(N5388) );
  CMXI2X1 U19980 ( .A0(n10106), .A1(n10100), .S(n4125), .Z(n10113) );
  CMX2X1 U19981 ( .A0(n10101), .A1(n10113), .S(n3773), .Z(n10126) );
  CMXI2X1 U19982 ( .A0(n10102), .A1(n10126), .S(n3426), .Z(N5389) );
  CMXI2X1 U19983 ( .A0(n10109), .A1(n10103), .S(n4125), .Z(n10116) );
  CMX2X1 U19984 ( .A0(n10104), .A1(n10116), .S(n3774), .Z(n10132) );
  CMXI2X1 U19985 ( .A0(n10105), .A1(n10132), .S(n3426), .Z(N5390) );
  CMXI2X1 U19986 ( .A0(n10112), .A1(n10106), .S(n4125), .Z(n10119) );
  CMX2X1 U19987 ( .A0(n10107), .A1(n10119), .S(n3775), .Z(n10135) );
  CMXI2X1 U19988 ( .A0(n10108), .A1(n10135), .S(n3425), .Z(N5391) );
  CMXI2X1 U19989 ( .A0(n10115), .A1(n10109), .S(n4125), .Z(n10122) );
  CMX2X1 U19990 ( .A0(n10110), .A1(n10122), .S(n3776), .Z(n10138) );
  CMXI2X1 U19991 ( .A0(n10111), .A1(n10138), .S(n3425), .Z(N5392) );
  CMXI2X1 U19992 ( .A0(n10118), .A1(n10112), .S(n4125), .Z(n10125) );
  CMX2X1 U19993 ( .A0(n10113), .A1(n10125), .S(n3777), .Z(n10141) );
  CMXI2X1 U19994 ( .A0(n10114), .A1(n10141), .S(n3425), .Z(N5393) );
  CMXI2X1 U19995 ( .A0(n10121), .A1(n10115), .S(n4125), .Z(n10131) );
  CMX2X1 U19996 ( .A0(n10116), .A1(n10131), .S(n3790), .Z(n10144) );
  CMXI2X1 U19997 ( .A0(n10117), .A1(n10144), .S(n3425), .Z(N5394) );
  CMXI2X1 U19998 ( .A0(n10124), .A1(n10118), .S(n4125), .Z(n10134) );
  CMX2X1 U19999 ( .A0(n10119), .A1(n10134), .S(n3791), .Z(n10147) );
  CMXI2X1 U20000 ( .A0(n10120), .A1(n10147), .S(n3425), .Z(N5395) );
  CMXI2X1 U20001 ( .A0(n10130), .A1(n10121), .S(n4125), .Z(n10137) );
  CMX2X1 U20002 ( .A0(n10122), .A1(n10137), .S(n3792), .Z(n10150) );
  CMXI2X1 U20003 ( .A0(n10123), .A1(n10150), .S(n3425), .Z(N5396) );
  CMXI2X1 U20004 ( .A0(n10133), .A1(n10124), .S(n4125), .Z(n10140) );
  CMX2X1 U20005 ( .A0(n10125), .A1(n10140), .S(n3793), .Z(n10153) );
  CMXI2X1 U20006 ( .A0(n10126), .A1(n10153), .S(n3428), .Z(N5397) );
  CMX2X1 U20007 ( .A0(N8242), .A1(N8241), .S(n4243), .Z(n10193) );
  CMXI2X1 U20008 ( .A0(n10193), .A1(n10127), .S(n4125), .Z(n10260) );
  CMX2X1 U20009 ( .A0(n10128), .A1(n10260), .S(n3794), .Z(n10400) );
  CMXI2X1 U20010 ( .A0(n10129), .A1(n10400), .S(n3428), .Z(N5181) );
  CMXI2X1 U20011 ( .A0(n10136), .A1(n10130), .S(n4125), .Z(n10143) );
  CMX2X1 U20012 ( .A0(n10131), .A1(n10143), .S(n3795), .Z(n10156) );
  CMXI2X1 U20013 ( .A0(n10132), .A1(n10156), .S(n3428), .Z(N5398) );
  CMXI2X1 U20014 ( .A0(n10139), .A1(n10133), .S(n4125), .Z(n10146) );
  CMX2X1 U20015 ( .A0(n10134), .A1(n10146), .S(n3796), .Z(n10159) );
  CMXI2X1 U20016 ( .A0(n10135), .A1(n10159), .S(n3428), .Z(N5399) );
  CMX2X1 U20017 ( .A0(N8023), .A1(N8022), .S(n4242), .Z(n10142) );
  CMXI2X1 U20018 ( .A0(n10142), .A1(n10136), .S(n4125), .Z(n10149) );
  CMX2X1 U20019 ( .A0(n10137), .A1(n10149), .S(n3797), .Z(n10165) );
  CMXI2X1 U20020 ( .A0(n10138), .A1(n10165), .S(n3428), .Z(N5400) );
  CMX2X1 U20021 ( .A0(N8022), .A1(N8021), .S(n4242), .Z(n10145) );
  CMXI2X1 U20022 ( .A0(n10145), .A1(n10139), .S(n4125), .Z(n10152) );
  CMX2X1 U20023 ( .A0(n10140), .A1(n10152), .S(n3805), .Z(n10168) );
  CMXI2X1 U20024 ( .A0(n10141), .A1(n10168), .S(n3428), .Z(N5401) );
  CMX2X1 U20025 ( .A0(N8021), .A1(N8020), .S(n4242), .Z(n10148) );
  CMXI2X1 U20026 ( .A0(n10148), .A1(n10142), .S(n4125), .Z(n10155) );
  CMX2X1 U20027 ( .A0(n10143), .A1(n10155), .S(n3806), .Z(n10171) );
  CMXI2X1 U20028 ( .A0(n10144), .A1(n10171), .S(n3428), .Z(N5402) );
  CMX2X1 U20029 ( .A0(N8020), .A1(N8019), .S(n4242), .Z(n10151) );
  CMXI2X1 U20030 ( .A0(n10151), .A1(n10145), .S(n4125), .Z(n10158) );
  CMX2X1 U20031 ( .A0(n10146), .A1(n10158), .S(n3790), .Z(n10174) );
  CMXI2X1 U20032 ( .A0(n10147), .A1(n10174), .S(n3428), .Z(N5403) );
  CMXI2X1 U20033 ( .A0(n10154), .A1(n10148), .S(n4124), .Z(n10164) );
  CMX2X1 U20034 ( .A0(n10149), .A1(n10164), .S(n3791), .Z(n10177) );
  CMXI2X1 U20035 ( .A0(n10150), .A1(n10177), .S(n3427), .Z(N5404) );
  CMXI2X1 U20036 ( .A0(n10157), .A1(n10151), .S(n4124), .Z(n10167) );
  CMX2X1 U20037 ( .A0(n10152), .A1(n10167), .S(n3773), .Z(n10180) );
  CMXI2X1 U20038 ( .A0(n10153), .A1(n10180), .S(n3427), .Z(N5405) );
  CMXI2X1 U20039 ( .A0(n10163), .A1(n10154), .S(n4124), .Z(n10170) );
  CMX2X1 U20040 ( .A0(n10155), .A1(n10170), .S(n3774), .Z(n10183) );
  CMXI2X1 U20041 ( .A0(n10156), .A1(n10183), .S(n3427), .Z(N5406) );
  CMXI2X1 U20042 ( .A0(n10166), .A1(n10157), .S(n4124), .Z(n10173) );
  CMX2X1 U20043 ( .A0(n10158), .A1(n10173), .S(n3775), .Z(n10186) );
  CMXI2X1 U20044 ( .A0(n10159), .A1(n10186), .S(n3427), .Z(N5407) );
  CMX2X1 U20045 ( .A0(N8241), .A1(N8240), .S(n4242), .Z(n10226) );
  CMXI2X1 U20046 ( .A0(n10226), .A1(n10160), .S(n4124), .Z(n10293) );
  CMX2X1 U20047 ( .A0(n10161), .A1(n10293), .S(n3776), .Z(n10433) );
  CMXI2X1 U20048 ( .A0(n10162), .A1(n10433), .S(n3427), .Z(N5182) );
  CMX2X1 U20049 ( .A0(N8015), .A1(N8014), .S(n4252), .Z(n10169) );
  CMXI2X1 U20050 ( .A0(n10169), .A1(n10163), .S(n4124), .Z(n10176) );
  CMX2X1 U20051 ( .A0(n10164), .A1(n10176), .S(n3777), .Z(n10189) );
  CMXI2X1 U20052 ( .A0(n10165), .A1(n10189), .S(n3427), .Z(N5408) );
  CMX2X1 U20053 ( .A0(N8014), .A1(N8013), .S(n4247), .Z(n10172) );
  CMXI2X1 U20054 ( .A0(n10172), .A1(n10166), .S(n4124), .Z(n10179) );
  CMX2X1 U20055 ( .A0(n10167), .A1(n10179), .S(n3811), .Z(n10192) );
  CMXI2X1 U20056 ( .A0(n10168), .A1(n10192), .S(n3427), .Z(N5409) );
  CMXI2X1 U20057 ( .A0(n10175), .A1(n10169), .S(n4124), .Z(n10182) );
  CMX2X1 U20058 ( .A0(n10170), .A1(n10182), .S(n3807), .Z(n10198) );
  CMXI2X1 U20059 ( .A0(n10171), .A1(n10198), .S(n3427), .Z(N5410) );
  CMXI2X1 U20060 ( .A0(n10178), .A1(n10172), .S(n4124), .Z(n10185) );
  CMX2X1 U20061 ( .A0(n10173), .A1(n10185), .S(n3808), .Z(n10201) );
  CMXI2X1 U20062 ( .A0(n10174), .A1(n10201), .S(n3427), .Z(N5411) );
  CMXI2X1 U20063 ( .A0(n10181), .A1(n10175), .S(n4124), .Z(n10188) );
  CMX2X1 U20064 ( .A0(n10176), .A1(n10188), .S(n3809), .Z(n10204) );
  CMXI2X1 U20065 ( .A0(n10177), .A1(n10204), .S(n3427), .Z(N5412) );
  CMXI2X1 U20066 ( .A0(n10184), .A1(n10178), .S(n4124), .Z(n10191) );
  CMX2X1 U20067 ( .A0(n10179), .A1(n10191), .S(n3810), .Z(n10207) );
  CMXI2X1 U20068 ( .A0(n10180), .A1(n10207), .S(n3395), .Z(N5413) );
  CMX2X1 U20069 ( .A0(N8009), .A1(N8008), .S(n4253), .Z(n10187) );
  CMXI2X1 U20070 ( .A0(n10187), .A1(n10181), .S(n4124), .Z(n10197) );
  CMX2X1 U20071 ( .A0(n10182), .A1(n10197), .S(n3811), .Z(n10210) );
  CMXI2X1 U20072 ( .A0(n10183), .A1(n10210), .S(n3395), .Z(N5414) );
  CMXI2X1 U20073 ( .A0(n10190), .A1(n10184), .S(n4124), .Z(n10200) );
  CMX2X1 U20074 ( .A0(n10185), .A1(n10200), .S(n3812), .Z(n10213) );
  CMXI2X1 U20075 ( .A0(n10186), .A1(n10213), .S(n3395), .Z(N5415) );
  CMX2X1 U20076 ( .A0(N8007), .A1(N8006), .S(n4230), .Z(n10196) );
  CMXI2X1 U20077 ( .A0(n10196), .A1(n10187), .S(n4124), .Z(n10203) );
  CMX2X1 U20078 ( .A0(n10188), .A1(n10203), .S(n4335), .Z(n10216) );
  CMXI2X1 U20079 ( .A0(n10189), .A1(n10216), .S(n3395), .Z(N5416) );
  CMX2X1 U20080 ( .A0(N8006), .A1(N8005), .S(n4247), .Z(n10199) );
  CMXI2X1 U20081 ( .A0(n10199), .A1(n10190), .S(n4124), .Z(n10206) );
  CMX2X1 U20082 ( .A0(n10191), .A1(n10206), .S(n3771), .Z(n10219) );
  CMXI2X1 U20083 ( .A0(n10192), .A1(n10219), .S(n3395), .Z(N5417) );
  CMX2X1 U20084 ( .A0(N8240), .A1(N8239), .S(n4241), .Z(n10259) );
  CMXI2X1 U20085 ( .A0(n10259), .A1(n10193), .S(n4124), .Z(n10326) );
  CMX2X1 U20086 ( .A0(n10194), .A1(n10326), .S(n3772), .Z(n10466) );
  CMXI2X1 U20087 ( .A0(n10195), .A1(n10466), .S(n3395), .Z(N5183) );
  CMXI2X1 U20088 ( .A0(n10202), .A1(n10196), .S(n4123), .Z(n10209) );
  CMX2X1 U20089 ( .A0(n10197), .A1(n10209), .S(n3773), .Z(n10222) );
  CMXI2X1 U20090 ( .A0(n10198), .A1(n10222), .S(n3395), .Z(N5418) );
  CMXI2X1 U20091 ( .A0(n10205), .A1(n10199), .S(n4123), .Z(n10212) );
  CMX2X1 U20092 ( .A0(n10200), .A1(n10212), .S(n3774), .Z(n10225) );
  CMXI2X1 U20093 ( .A0(n10201), .A1(n10225), .S(n3395), .Z(N5419) );
  CMX2X1 U20094 ( .A0(N8003), .A1(N8002), .S(n4241), .Z(n10208) );
  CMXI2X1 U20095 ( .A0(n10208), .A1(n10202), .S(n4123), .Z(n10215) );
  CMX2X1 U20096 ( .A0(n10203), .A1(n10215), .S(n3775), .Z(n10231) );
  CMXI2X1 U20097 ( .A0(n10204), .A1(n10231), .S(n3395), .Z(N5420) );
  CMX2X1 U20098 ( .A0(N8002), .A1(N8001), .S(n4241), .Z(n10211) );
  CMXI2X1 U20099 ( .A0(n10211), .A1(n10205), .S(n4123), .Z(n10218) );
  CMX2X1 U20100 ( .A0(n10206), .A1(n10218), .S(n3776), .Z(n10234) );
  CMXI2X1 U20101 ( .A0(n10207), .A1(n10234), .S(n3394), .Z(N5421) );
  CMX2X1 U20102 ( .A0(N8001), .A1(N8000), .S(n4241), .Z(n10214) );
  CMXI2X1 U20103 ( .A0(n10214), .A1(n10208), .S(n4123), .Z(n10221) );
  CMX2X1 U20104 ( .A0(n10209), .A1(n10221), .S(n3777), .Z(n10237) );
  CMXI2X1 U20105 ( .A0(n10210), .A1(n10237), .S(n3394), .Z(N5422) );
  CMX2X1 U20106 ( .A0(N8000), .A1(N7999), .S(n4241), .Z(n10217) );
  CMXI2X1 U20107 ( .A0(n10217), .A1(n10211), .S(n4123), .Z(n10224) );
  CMX2X1 U20108 ( .A0(n10212), .A1(n10224), .S(n3790), .Z(n10240) );
  CMXI2X1 U20109 ( .A0(n10213), .A1(n10240), .S(n3394), .Z(N5423) );
  CMX2X1 U20110 ( .A0(N7999), .A1(N7998), .S(n4241), .Z(n10220) );
  CMXI2X1 U20111 ( .A0(n10220), .A1(n10214), .S(n4123), .Z(n10230) );
  CMX2X1 U20112 ( .A0(n10215), .A1(n10230), .S(n3791), .Z(n10243) );
  CMXI2X1 U20113 ( .A0(n10216), .A1(n10243), .S(n3403), .Z(N5424) );
  CMX2X1 U20114 ( .A0(N7998), .A1(N7997), .S(n4241), .Z(n10223) );
  CMXI2X1 U20115 ( .A0(n10223), .A1(n10217), .S(n4123), .Z(n10233) );
  CMX2X1 U20116 ( .A0(n10218), .A1(n10233), .S(n3792), .Z(n10246) );
  CMXI2X1 U20117 ( .A0(n10219), .A1(n10246), .S(n3429), .Z(N5425) );
  CMX2X1 U20118 ( .A0(N7997), .A1(N7996), .S(n4241), .Z(n10229) );
  CMXI2X1 U20119 ( .A0(n10229), .A1(n10220), .S(n4123), .Z(n10236) );
  CMX2X1 U20120 ( .A0(n10221), .A1(n10236), .S(n3790), .Z(n10249) );
  CMXI2X1 U20121 ( .A0(n10222), .A1(n10249), .S(n3429), .Z(N5426) );
  CMX2X1 U20122 ( .A0(N7996), .A1(N7995), .S(n4241), .Z(n10232) );
  CMXI2X1 U20123 ( .A0(n10232), .A1(n10223), .S(n4123), .Z(n10239) );
  CMX2X1 U20124 ( .A0(n10224), .A1(n10239), .S(n3791), .Z(n10252) );
  CMXI2X1 U20125 ( .A0(n10225), .A1(n10252), .S(n3428), .Z(N5427) );
  CMX2X1 U20126 ( .A0(N8239), .A1(N8238), .S(n4243), .Z(n10292) );
  CMXI2X1 U20127 ( .A0(n10292), .A1(n10226), .S(n4123), .Z(n10366) );
  CMX2X1 U20128 ( .A0(n10227), .A1(n10366), .S(n3792), .Z(n10499) );
  CMXI2X1 U20129 ( .A0(n10228), .A1(n10499), .S(n3428), .Z(N5184) );
  CMXI2X1 U20130 ( .A0(n10235), .A1(n10229), .S(n4123), .Z(n10242) );
  CMX2X1 U20131 ( .A0(n10230), .A1(n10242), .S(n3793), .Z(n10255) );
  CMXI2X1 U20132 ( .A0(n10231), .A1(n10255), .S(n3428), .Z(N5428) );
  CMXI2X1 U20133 ( .A0(n10238), .A1(n10232), .S(n4123), .Z(n10245) );
  CMX2X1 U20134 ( .A0(n10233), .A1(n10245), .S(n3794), .Z(n10258) );
  CMXI2X1 U20135 ( .A0(n10234), .A1(n10258), .S(n3397), .Z(N5429) );
  CMX2X1 U20136 ( .A0(N7993), .A1(N7992), .S(n4245), .Z(n10241) );
  CMXI2X1 U20137 ( .A0(n10241), .A1(n10235), .S(n4123), .Z(n10248) );
  CMX2X1 U20138 ( .A0(n10236), .A1(n10248), .S(n3812), .Z(n10264) );
  CMXI2X1 U20139 ( .A0(n10237), .A1(n10264), .S(n3397), .Z(N5430) );
  CMX2X1 U20140 ( .A0(N7992), .A1(N7991), .S(n4244), .Z(n10244) );
  CMXI2X1 U20141 ( .A0(n10244), .A1(n10238), .S(n4123), .Z(n10251) );
  CMX2X1 U20142 ( .A0(n10239), .A1(n10251), .S(n3792), .Z(n10267) );
  CMXI2X1 U20143 ( .A0(n10240), .A1(n10267), .S(n3397), .Z(N5431) );
  CMXI2X1 U20144 ( .A0(n10247), .A1(n10241), .S(n4123), .Z(n10254) );
  CMX2X1 U20145 ( .A0(n10242), .A1(n10254), .S(n3793), .Z(n10270) );
  CMXI2X1 U20146 ( .A0(n10243), .A1(n10270), .S(n3397), .Z(N5432) );
  CMXI2X1 U20147 ( .A0(n10250), .A1(n10244), .S(n4122), .Z(n10257) );
  CMX2X1 U20148 ( .A0(n10245), .A1(n10257), .S(n3794), .Z(n10273) );
  CMXI2X1 U20149 ( .A0(n10246), .A1(n10273), .S(n3397), .Z(N5433) );
  CMXI2X1 U20150 ( .A0(n10253), .A1(n10247), .S(n4122), .Z(n10263) );
  CMX2X1 U20151 ( .A0(n10248), .A1(n10263), .S(n3795), .Z(n10276) );
  CMXI2X1 U20152 ( .A0(n10249), .A1(n10276), .S(n3396), .Z(N5434) );
  CMXI2X1 U20153 ( .A0(n10256), .A1(n10250), .S(n4122), .Z(n10266) );
  CMX2X1 U20154 ( .A0(n10251), .A1(n10266), .S(n3796), .Z(n10279) );
  CMXI2X1 U20155 ( .A0(n10252), .A1(n10279), .S(n3396), .Z(N5435) );
  CMXI2X1 U20156 ( .A0(n10262), .A1(n10253), .S(n4122), .Z(n10269) );
  CMX2X1 U20157 ( .A0(n10254), .A1(n10269), .S(n3797), .Z(n10282) );
  CMXI2X1 U20158 ( .A0(n10255), .A1(n10282), .S(n3396), .Z(N5436) );
  CMXI2X1 U20159 ( .A0(n10265), .A1(n10256), .S(n4122), .Z(n10272) );
  CMX2X1 U20160 ( .A0(n10257), .A1(n10272), .S(n3805), .Z(n10285) );
  CMXI2X1 U20161 ( .A0(n10258), .A1(n10285), .S(n3396), .Z(N5437) );
  CMX2X1 U20162 ( .A0(N8238), .A1(N8237), .S(n4240), .Z(n10325) );
  CMXI2X1 U20163 ( .A0(n10325), .A1(n10259), .S(n4122), .Z(n10399) );
  CMX2X1 U20164 ( .A0(n10260), .A1(n10399), .S(n3806), .Z(n10532) );
  CMXI2X1 U20165 ( .A0(n10261), .A1(n10532), .S(n3396), .Z(N5185) );
  CMXI2X1 U20166 ( .A0(n10268), .A1(n10262), .S(n4122), .Z(n10275) );
  CMX2X1 U20167 ( .A0(n10263), .A1(n10275), .S(n3807), .Z(n10288) );
  CMXI2X1 U20168 ( .A0(n10264), .A1(n10288), .S(n3396), .Z(N5438) );
  CMXI2X1 U20169 ( .A0(n10271), .A1(n10265), .S(n4122), .Z(n10278) );
  CMX2X1 U20170 ( .A0(n10266), .A1(n10278), .S(n3808), .Z(n10291) );
  CMXI2X1 U20171 ( .A0(n10267), .A1(n10291), .S(n3396), .Z(N5439) );
  CMXI2X1 U20172 ( .A0(n10274), .A1(n10268), .S(n4122), .Z(n10281) );
  CMX2X1 U20173 ( .A0(n10269), .A1(n10281), .S(n3809), .Z(n10297) );
  CMXI2X1 U20174 ( .A0(n10270), .A1(n10297), .S(n3396), .Z(N5440) );
  CMXI2X1 U20175 ( .A0(n10277), .A1(n10271), .S(n4122), .Z(n10284) );
  CMX2X1 U20176 ( .A0(n10272), .A1(n10284), .S(n3810), .Z(n10300) );
  CMXI2X1 U20177 ( .A0(n10273), .A1(n10300), .S(n3396), .Z(N5441) );
  CMXI2X1 U20178 ( .A0(n10280), .A1(n10274), .S(n4122), .Z(n10287) );
  CMX2X1 U20179 ( .A0(n10275), .A1(n10287), .S(n3811), .Z(n10303) );
  CMXI2X1 U20180 ( .A0(n10276), .A1(n10303), .S(n3396), .Z(N5442) );
  CMXI2X1 U20181 ( .A0(n10283), .A1(n10277), .S(n4122), .Z(n10290) );
  CMX2X1 U20182 ( .A0(n10278), .A1(n10290), .S(n3812), .Z(n10306) );
  CMXI2X1 U20183 ( .A0(n10279), .A1(n10306), .S(n3395), .Z(N5443) );
  CMXI2X1 U20184 ( .A0(n10286), .A1(n10280), .S(n4122), .Z(n10296) );
  CMX2X1 U20185 ( .A0(n10281), .A1(n10296), .S(n4334), .Z(n10309) );
  CMXI2X1 U20186 ( .A0(n10282), .A1(n10309), .S(n3395), .Z(N5444) );
  CMXI2X1 U20187 ( .A0(n10289), .A1(n10283), .S(n4122), .Z(n10299) );
  CMX2X1 U20188 ( .A0(n10284), .A1(n10299), .S(n3771), .Z(n10312) );
  CMXI2X1 U20189 ( .A0(n10285), .A1(n10312), .S(n3399), .Z(N5445) );
  CMXI2X1 U20190 ( .A0(n10295), .A1(n10286), .S(n4122), .Z(n10302) );
  CMX2X1 U20191 ( .A0(n10287), .A1(n10302), .S(n3792), .Z(n10315) );
  CMXI2X1 U20192 ( .A0(n10288), .A1(n10315), .S(n3398), .Z(N5446) );
  CMXI2X1 U20193 ( .A0(n10298), .A1(n10289), .S(n4122), .Z(n10305) );
  CMX2X1 U20194 ( .A0(n10290), .A1(n10305), .S(n3793), .Z(n10318) );
  CMXI2X1 U20195 ( .A0(n10291), .A1(n10318), .S(n3398), .Z(N5447) );
  CMX2X1 U20196 ( .A0(N8237), .A1(N8236), .S(n4239), .Z(n10365) );
  CMXI2X1 U20197 ( .A0(n10365), .A1(n10292), .S(n4121), .Z(n10432) );
  CMX2X1 U20198 ( .A0(n10293), .A1(n10432), .S(n3795), .Z(n10565) );
  CMXI2X1 U20199 ( .A0(n10294), .A1(n10565), .S(n3398), .Z(N5186) );
  CMXI2X1 U20200 ( .A0(n10301), .A1(n10295), .S(n4121), .Z(n10308) );
  CMX2X1 U20201 ( .A0(n10296), .A1(n10308), .S(n3796), .Z(n10321) );
  CMXI2X1 U20202 ( .A0(n10297), .A1(n10321), .S(n3398), .Z(N5448) );
  CMXI2X1 U20203 ( .A0(n10304), .A1(n10298), .S(n4121), .Z(n10311) );
  CMX2X1 U20204 ( .A0(n10299), .A1(n10311), .S(n3797), .Z(n10324) );
  CMXI2X1 U20205 ( .A0(n10300), .A1(n10324), .S(n3398), .Z(N5449) );
  CMXI2X1 U20206 ( .A0(n10307), .A1(n10301), .S(n4121), .Z(n10314) );
  CMX2X1 U20207 ( .A0(n10302), .A1(n10314), .S(n3805), .Z(n10337) );
  CMXI2X1 U20208 ( .A0(n10303), .A1(n10337), .S(n3398), .Z(N5450) );
  CMXI2X1 U20209 ( .A0(n10310), .A1(n10304), .S(n4121), .Z(n10317) );
  CMX2X1 U20210 ( .A0(n10305), .A1(n10317), .S(n3806), .Z(n10340) );
  CMXI2X1 U20211 ( .A0(n10306), .A1(n10340), .S(n3398), .Z(N5451) );
  CMXI2X1 U20212 ( .A0(n10313), .A1(n10307), .S(n4121), .Z(n10320) );
  CMX2X1 U20213 ( .A0(n10308), .A1(n10320), .S(n4312), .Z(n10343) );
  CMXI2X1 U20214 ( .A0(n10309), .A1(n10343), .S(n3398), .Z(N5452) );
  CMXI2X1 U20215 ( .A0(n10316), .A1(n10310), .S(n4121), .Z(n10323) );
  CMX2X1 U20216 ( .A0(n10311), .A1(n10323), .S(n3772), .Z(n10346) );
  CMXI2X1 U20217 ( .A0(n10312), .A1(n10346), .S(n3398), .Z(N5453) );
  CMX2X1 U20218 ( .A0(N7969), .A1(N7968), .S(n4239), .Z(n10319) );
  CMXI2X1 U20219 ( .A0(n10319), .A1(n10313), .S(n4121), .Z(n10336) );
  CMX2X1 U20220 ( .A0(n10314), .A1(n10336), .S(n3773), .Z(n10349) );
  CMXI2X1 U20221 ( .A0(n10315), .A1(n10349), .S(n3398), .Z(N5454) );
  CMXI2X1 U20222 ( .A0(n10322), .A1(n10316), .S(n4121), .Z(n10339) );
  CMX2X1 U20223 ( .A0(n10317), .A1(n10339), .S(n3774), .Z(n10352) );
  CMXI2X1 U20224 ( .A0(n10318), .A1(n10352), .S(n3398), .Z(N5455) );
  CMXI2X1 U20225 ( .A0(n10335), .A1(n10319), .S(n4121), .Z(n10342) );
  CMX2X1 U20226 ( .A0(n10320), .A1(n10342), .S(n3775), .Z(n10355) );
  CMXI2X1 U20227 ( .A0(n10321), .A1(n10355), .S(n3397), .Z(N5456) );
  CMXI2X1 U20228 ( .A0(n10338), .A1(n10322), .S(n4121), .Z(n10345) );
  CMX2X1 U20229 ( .A0(n10323), .A1(n10345), .S(n3776), .Z(n10358) );
  CMXI2X1 U20230 ( .A0(n10324), .A1(n10358), .S(n3397), .Z(N5457) );
  CMX2X1 U20231 ( .A0(N8236), .A1(N8235), .S(n4255), .Z(n10398) );
  CMXI2X1 U20232 ( .A0(n10398), .A1(n10325), .S(n4121), .Z(n10465) );
  CMX2X1 U20233 ( .A0(n10326), .A1(n10465), .S(n3777), .Z(n10598) );
  CMXI2X1 U20234 ( .A0(n10327), .A1(n10598), .S(n3397), .Z(N5187) );
  CMXI2X1 U20235 ( .A0(n10329), .A1(n10328), .S(n4121), .Z(n11671) );
  CMXI2X1 U20236 ( .A0(n10331), .A1(n10330), .S(n4121), .Z(n10332) );
  CMXI2X1 U20237 ( .A0(n11671), .A1(n10332), .S(n3798), .Z(n10334) );
  CMXI2X1 U20238 ( .A0(n10334), .A1(n10333), .S(n3397), .Z(N5160) );
  CMXI2X1 U20239 ( .A0(n10341), .A1(n10335), .S(n4121), .Z(n10348) );
  CMX2X1 U20240 ( .A0(n10336), .A1(n10348), .S(n3790), .Z(n10361) );
  CMXI2X1 U20241 ( .A0(n10337), .A1(n10361), .S(n3397), .Z(N5458) );
  CMXI2X1 U20242 ( .A0(n10344), .A1(n10338), .S(n4121), .Z(n10351) );
  CMX2X1 U20243 ( .A0(n10339), .A1(n10351), .S(n3791), .Z(n10364) );
  CMXI2X1 U20244 ( .A0(n10340), .A1(n10364), .S(n3397), .Z(N5459) );
  CMXI2X1 U20245 ( .A0(n10347), .A1(n10341), .S(n4120), .Z(n10354) );
  CMX2X1 U20246 ( .A0(n10342), .A1(n10354), .S(n3792), .Z(n10370) );
  CMXI2X1 U20247 ( .A0(n10343), .A1(n10370), .S(n3400), .Z(N5460) );
  CMXI2X1 U20248 ( .A0(n10350), .A1(n10344), .S(n4120), .Z(n10357) );
  CMX2X1 U20249 ( .A0(n10345), .A1(n10357), .S(n3793), .Z(n10373) );
  CMXI2X1 U20250 ( .A0(n10346), .A1(n10373), .S(n3400), .Z(N5461) );
  CMXI2X1 U20251 ( .A0(n10353), .A1(n10347), .S(n4120), .Z(n10360) );
  CMX2X1 U20252 ( .A0(n10348), .A1(n10360), .S(n3794), .Z(n10376) );
  CMXI2X1 U20253 ( .A0(n10349), .A1(n10376), .S(n3400), .Z(N5462) );
  CMXI2X1 U20254 ( .A0(n10356), .A1(n10350), .S(n4120), .Z(n10363) );
  CMX2X1 U20255 ( .A0(n10351), .A1(n10363), .S(n3795), .Z(n10379) );
  CMXI2X1 U20256 ( .A0(n10352), .A1(n10379), .S(n3400), .Z(N5463) );
  CMX2X1 U20257 ( .A0(N7959), .A1(N7958), .S(n4250), .Z(n10359) );
  CMXI2X1 U20258 ( .A0(n10359), .A1(n10353), .S(n4120), .Z(n10369) );
  CMX2X1 U20259 ( .A0(n10354), .A1(n10369), .S(n3796), .Z(n10382) );
  CMXI2X1 U20260 ( .A0(n10355), .A1(n10382), .S(n3400), .Z(N5464) );
  CMX2X1 U20261 ( .A0(N7958), .A1(N7957), .S(n4251), .Z(n10362) );
  CMXI2X1 U20262 ( .A0(n10362), .A1(n10356), .S(n4120), .Z(n10372) );
  CMX2X1 U20263 ( .A0(n10357), .A1(n10372), .S(n3797), .Z(n10385) );
  CMXI2X1 U20264 ( .A0(n10358), .A1(n10385), .S(n3400), .Z(N5465) );
  CMX2X1 U20265 ( .A0(N7957), .A1(N7956), .S(n4249), .Z(n10368) );
  CMXI2X1 U20266 ( .A0(n10368), .A1(n10359), .S(n4120), .Z(n10375) );
  CMX2X1 U20267 ( .A0(n10360), .A1(n10375), .S(n3805), .Z(n10388) );
  CMXI2X1 U20268 ( .A0(n10361), .A1(n10388), .S(n3400), .Z(N5466) );
  CMX2X1 U20269 ( .A0(N7956), .A1(N7955), .S(n4280), .Z(n10371) );
  CMXI2X1 U20270 ( .A0(n10371), .A1(n10362), .S(n4120), .Z(n10378) );
  CMX2X1 U20271 ( .A0(n10363), .A1(n10378), .S(n3806), .Z(n10391) );
  CMXI2X1 U20272 ( .A0(n10364), .A1(n10391), .S(n3400), .Z(N5467) );
  CMX2X1 U20273 ( .A0(N8235), .A1(N8234), .S(n4248), .Z(n10431) );
  CMXI2X1 U20274 ( .A0(n10431), .A1(n10365), .S(n4120), .Z(n10498) );
  CMX2X1 U20275 ( .A0(n10366), .A1(n10498), .S(n3793), .Z(n10631) );
  CMXI2X1 U20276 ( .A0(n10367), .A1(n10631), .S(n3399), .Z(N5188) );
  CMXI2X1 U20277 ( .A0(n10374), .A1(n10368), .S(n4120), .Z(n10381) );
  CMX2X1 U20278 ( .A0(n10369), .A1(n10381), .S(n3794), .Z(n10394) );
  CMXI2X1 U20279 ( .A0(n10370), .A1(n10394), .S(n3399), .Z(N5468) );
  CMXI2X1 U20280 ( .A0(n10377), .A1(n10371), .S(n4120), .Z(n10384) );
  CMX2X1 U20281 ( .A0(n10372), .A1(n10384), .S(n3807), .Z(n10397) );
  CMXI2X1 U20282 ( .A0(n10373), .A1(n10397), .S(n3399), .Z(N5469) );
  CMXI2X1 U20283 ( .A0(n10380), .A1(n10374), .S(n4120), .Z(n10387) );
  CMX2X1 U20284 ( .A0(n10375), .A1(n10387), .S(n3808), .Z(n10403) );
  CMXI2X1 U20285 ( .A0(n10376), .A1(n10403), .S(n3399), .Z(N5470) );
  CMXI2X1 U20286 ( .A0(n10383), .A1(n10377), .S(n4120), .Z(n10390) );
  CMX2X1 U20287 ( .A0(n10378), .A1(n10390), .S(n3771), .Z(n10406) );
  CMXI2X1 U20288 ( .A0(n10379), .A1(n10406), .S(n3399), .Z(N5471) );
  CMX2X1 U20289 ( .A0(N7951), .A1(N7950), .S(n4248), .Z(n10386) );
  CMXI2X1 U20290 ( .A0(n10386), .A1(n10380), .S(n4120), .Z(n10393) );
  CMX2X1 U20291 ( .A0(n10381), .A1(n10393), .S(n3812), .Z(n10409) );
  CMXI2X1 U20292 ( .A0(n10382), .A1(n10409), .S(n3399), .Z(N5472) );
  CMX2X1 U20293 ( .A0(N7950), .A1(N7949), .S(n4233), .Z(n10389) );
  CMXI2X1 U20294 ( .A0(n10389), .A1(n10383), .S(n4120), .Z(n10396) );
  CMX2X1 U20295 ( .A0(n10384), .A1(n10396), .S(n3805), .Z(n10412) );
  CMXI2X1 U20296 ( .A0(n10385), .A1(n10412), .S(n3399), .Z(N5473) );
  CMXI2X1 U20297 ( .A0(n10392), .A1(n10386), .S(n4120), .Z(n10402) );
  CMX2X1 U20298 ( .A0(n10387), .A1(n10402), .S(n4309), .Z(n10415) );
  CMXI2X1 U20299 ( .A0(n10388), .A1(n10415), .S(n3399), .Z(N5474) );
  CMXI2X1 U20300 ( .A0(n10395), .A1(n10389), .S(n4119), .Z(n10405) );
  CMX2X1 U20301 ( .A0(n10390), .A1(n10405), .S(n3771), .Z(n10418) );
  CMXI2X1 U20302 ( .A0(n10391), .A1(n10418), .S(n3399), .Z(N5475) );
  CMX2X1 U20303 ( .A0(N7947), .A1(N7946), .S(n4231), .Z(n10401) );
  CMXI2X1 U20304 ( .A0(n10401), .A1(n10392), .S(n4119), .Z(n10408) );
  CMX2X1 U20305 ( .A0(n10393), .A1(n10408), .S(n3772), .Z(n10421) );
  CMXI2X1 U20306 ( .A0(n10394), .A1(n10421), .S(n3399), .Z(N5476) );
  CMX2X1 U20307 ( .A0(N7946), .A1(N7945), .S(n4232), .Z(n10404) );
  CMXI2X1 U20308 ( .A0(n10404), .A1(n10395), .S(n4119), .Z(n10411) );
  CMX2X1 U20309 ( .A0(n10396), .A1(n10411), .S(n3773), .Z(n10424) );
  CMXI2X1 U20310 ( .A0(n10397), .A1(n10424), .S(n3402), .Z(N5477) );
  CMX2X1 U20311 ( .A0(N8234), .A1(N8233), .S(n4238), .Z(n10464) );
  CMXI2X1 U20312 ( .A0(n10464), .A1(n10398), .S(n4119), .Z(n10531) );
  CMX2X1 U20313 ( .A0(n10399), .A1(n10531), .S(n3774), .Z(n10664) );
  CMXI2X1 U20314 ( .A0(n10400), .A1(n10664), .S(n3402), .Z(N5189) );
  CMXI2X1 U20315 ( .A0(n10407), .A1(n10401), .S(n4119), .Z(n10414) );
  CMX2X1 U20316 ( .A0(n10402), .A1(n10414), .S(n3805), .Z(n10427) );
  CMXI2X1 U20317 ( .A0(n10403), .A1(n10427), .S(n3402), .Z(N5478) );
  CMXI2X1 U20318 ( .A0(n10410), .A1(n10404), .S(n4119), .Z(n10417) );
  CMX2X1 U20319 ( .A0(n10405), .A1(n10417), .S(n3772), .Z(n10430) );
  CMXI2X1 U20320 ( .A0(n10406), .A1(n10430), .S(n3402), .Z(N5479) );
  CMX2X1 U20321 ( .A0(N7943), .A1(N7942), .S(n4238), .Z(n10413) );
  CMXI2X1 U20322 ( .A0(n10413), .A1(n10407), .S(n4119), .Z(n10420) );
  CMX2X1 U20323 ( .A0(n10408), .A1(n10420), .S(n3773), .Z(n10436) );
  CMXI2X1 U20324 ( .A0(n10409), .A1(n10436), .S(n3401), .Z(N5480) );
  CMX2X1 U20325 ( .A0(N7942), .A1(N7941), .S(n4238), .Z(n10416) );
  CMXI2X1 U20326 ( .A0(n10416), .A1(n10410), .S(n4119), .Z(n10423) );
  CMX2X1 U20327 ( .A0(n10411), .A1(n10423), .S(n3774), .Z(n10439) );
  CMXI2X1 U20328 ( .A0(n10412), .A1(n10439), .S(n3401), .Z(N5481) );
  CMXI2X1 U20329 ( .A0(n10419), .A1(n10413), .S(n4119), .Z(n10426) );
  CMX2X1 U20330 ( .A0(n10414), .A1(n10426), .S(n3775), .Z(n10442) );
  CMXI2X1 U20331 ( .A0(n10415), .A1(n10442), .S(n3401), .Z(N5482) );
  CMXI2X1 U20332 ( .A0(n10422), .A1(n10416), .S(n4119), .Z(n10429) );
  CMX2X1 U20333 ( .A0(n10417), .A1(n10429), .S(n3776), .Z(n10445) );
  CMXI2X1 U20334 ( .A0(n10418), .A1(n10445), .S(n3401), .Z(N5483) );
  CMX2X1 U20335 ( .A0(N7939), .A1(N7938), .S(n4238), .Z(n10425) );
  CMXI2X1 U20336 ( .A0(n10425), .A1(n10419), .S(n4119), .Z(n10435) );
  CMX2X1 U20337 ( .A0(n10420), .A1(n10435), .S(n3777), .Z(n10448) );
  CMXI2X1 U20338 ( .A0(n10421), .A1(n10448), .S(n3401), .Z(N5484) );
  CMX2X1 U20339 ( .A0(N7938), .A1(N7937), .S(n4238), .Z(n10428) );
  CMXI2X1 U20340 ( .A0(n10428), .A1(n10422), .S(n4119), .Z(n10438) );
  CMX2X1 U20341 ( .A0(n10423), .A1(n10438), .S(n3790), .Z(n10451) );
  CMXI2X1 U20342 ( .A0(n10424), .A1(n10451), .S(n3401), .Z(N5485) );
  CMX2X1 U20343 ( .A0(N7937), .A1(N7936), .S(n4238), .Z(n10434) );
  CMXI2X1 U20344 ( .A0(n10434), .A1(n10425), .S(n4119), .Z(n10441) );
  CMX2X1 U20345 ( .A0(n10426), .A1(n10441), .S(n3791), .Z(n10454) );
  CMXI2X1 U20346 ( .A0(n10427), .A1(n10454), .S(n3401), .Z(N5486) );
  CMX2X1 U20347 ( .A0(N7936), .A1(N7935), .S(n4238), .Z(n10437) );
  CMXI2X1 U20348 ( .A0(n10437), .A1(n10428), .S(n4119), .Z(n10444) );
  CMX2X1 U20349 ( .A0(n10429), .A1(n10444), .S(n3792), .Z(n10457) );
  CMXI2X1 U20350 ( .A0(n10430), .A1(n10457), .S(n3401), .Z(N5487) );
  CMX2X1 U20351 ( .A0(N8233), .A1(N8232), .S(n4237), .Z(n10497) );
  CMXI2X1 U20352 ( .A0(n10497), .A1(n10431), .S(n4119), .Z(n10564) );
  CMX2X1 U20353 ( .A0(n10432), .A1(n10564), .S(n3793), .Z(n10704) );
  CMXI2X1 U20354 ( .A0(n10433), .A1(n10704), .S(n3401), .Z(N5190) );
  CMX2X1 U20355 ( .A0(N7935), .A1(N7934), .S(n4237), .Z(n10440) );
  CMXI2X1 U20356 ( .A0(n10440), .A1(n10434), .S(n4119), .Z(n10447) );
  CMX2X1 U20357 ( .A0(n10435), .A1(n10447), .S(n3794), .Z(n10460) );
  CMXI2X1 U20358 ( .A0(n10436), .A1(n10460), .S(n3401), .Z(N5488) );
  CMX2X1 U20359 ( .A0(N7934), .A1(N7933), .S(n4237), .Z(n10443) );
  CMXI2X1 U20360 ( .A0(n10443), .A1(n10437), .S(n4118), .Z(n10450) );
  CMX2X1 U20361 ( .A0(n10438), .A1(n10450), .S(n3795), .Z(n10463) );
  CMXI2X1 U20362 ( .A0(n10439), .A1(n10463), .S(n3401), .Z(N5489) );
  CMX2X1 U20363 ( .A0(N7933), .A1(N7932), .S(n4237), .Z(n10446) );
  CMXI2X1 U20364 ( .A0(n10446), .A1(n10440), .S(n4118), .Z(n10453) );
  CMX2X1 U20365 ( .A0(n10441), .A1(n10453), .S(n3796), .Z(n10469) );
  CMXI2X1 U20366 ( .A0(n10442), .A1(n10469), .S(n3400), .Z(N5490) );
  CMX2X1 U20367 ( .A0(N7932), .A1(N7931), .S(n4237), .Z(n10449) );
  CMXI2X1 U20368 ( .A0(n10449), .A1(n10443), .S(n4118), .Z(n10456) );
  CMX2X1 U20369 ( .A0(n10444), .A1(n10456), .S(n3808), .Z(n10472) );
  CMXI2X1 U20370 ( .A0(n10445), .A1(n10472), .S(n3400), .Z(N5491) );
  CMXI2X1 U20371 ( .A0(n10452), .A1(n10446), .S(n4118), .Z(n10459) );
  CMX2X1 U20372 ( .A0(n10447), .A1(n10459), .S(n3807), .Z(n10475) );
  CMXI2X1 U20373 ( .A0(n10448), .A1(n10475), .S(n3400), .Z(N5492) );
  CMXI2X1 U20374 ( .A0(n10455), .A1(n10449), .S(n4118), .Z(n10462) );
  CMX2X1 U20375 ( .A0(n10450), .A1(n10462), .S(n3808), .Z(n10478) );
  CMXI2X1 U20376 ( .A0(n10451), .A1(n10478), .S(n3404), .Z(N5493) );
  CMX2X1 U20377 ( .A0(N7929), .A1(N7928), .S(n4237), .Z(n10458) );
  CMXI2X1 U20378 ( .A0(n10458), .A1(n10452), .S(n4118), .Z(n10468) );
  CMX2X1 U20379 ( .A0(n10453), .A1(n10468), .S(n3809), .Z(n10481) );
  CMXI2X1 U20380 ( .A0(n10454), .A1(n10481), .S(n3403), .Z(N5494) );
  CMX2X1 U20381 ( .A0(N7928), .A1(N7927), .S(n4237), .Z(n10461) );
  CMXI2X1 U20382 ( .A0(n10461), .A1(n10455), .S(n4118), .Z(n10471) );
  CMX2X1 U20383 ( .A0(n10456), .A1(n10471), .S(n3810), .Z(n10484) );
  CMXI2X1 U20384 ( .A0(n10457), .A1(n10484), .S(n3403), .Z(N5495) );
  CMXI2X1 U20385 ( .A0(n10467), .A1(n10458), .S(n4118), .Z(n10474) );
  CMX2X1 U20386 ( .A0(n10459), .A1(n10474), .S(n3811), .Z(n10487) );
  CMXI2X1 U20387 ( .A0(n10460), .A1(n10487), .S(n3403), .Z(N5496) );
  CMXI2X1 U20388 ( .A0(n10470), .A1(n10461), .S(n4118), .Z(n10477) );
  CMX2X1 U20389 ( .A0(n10462), .A1(n10477), .S(n3812), .Z(n10490) );
  CMXI2X1 U20390 ( .A0(n10463), .A1(n10490), .S(n3403), .Z(N5497) );
  CMX2X1 U20391 ( .A0(N8232), .A1(N8231), .S(n4236), .Z(n10530) );
  CMXI2X1 U20392 ( .A0(n10530), .A1(n10464), .S(n4118), .Z(n10597) );
  CMX2X1 U20393 ( .A0(n10465), .A1(n10597), .S(n4337), .Z(n10737) );
  CMXI2X1 U20394 ( .A0(n10466), .A1(n10737), .S(n3403), .Z(N5191) );
  CMXI2X1 U20395 ( .A0(n10473), .A1(n10467), .S(n4118), .Z(n10480) );
  CMX2X1 U20396 ( .A0(n10468), .A1(n10480), .S(n3771), .Z(n10493) );
  CMXI2X1 U20397 ( .A0(n10469), .A1(n10493), .S(n3403), .Z(N5498) );
  CMXI2X1 U20398 ( .A0(n10476), .A1(n10470), .S(n4118), .Z(n10483) );
  CMX2X1 U20399 ( .A0(n10471), .A1(n10483), .S(n3772), .Z(n10496) );
  CMXI2X1 U20400 ( .A0(n10472), .A1(n10496), .S(n3403), .Z(N5499) );
  CMXI2X1 U20401 ( .A0(n10479), .A1(n10473), .S(n4118), .Z(n10486) );
  CMX2X1 U20402 ( .A0(n10474), .A1(n10486), .S(n3773), .Z(n10502) );
  CMXI2X1 U20403 ( .A0(n10475), .A1(n10502), .S(n3403), .Z(N5500) );
  CMXI2X1 U20404 ( .A0(n10482), .A1(n10476), .S(n4118), .Z(n10489) );
  CMX2X1 U20405 ( .A0(n10477), .A1(n10489), .S(n3774), .Z(n10505) );
  CMXI2X1 U20406 ( .A0(n10478), .A1(n10505), .S(n3403), .Z(N5501) );
  CMXI2X1 U20407 ( .A0(n10485), .A1(n10479), .S(n4118), .Z(n10492) );
  CMX2X1 U20408 ( .A0(n10480), .A1(n10492), .S(n3775), .Z(n10508) );
  CMXI2X1 U20409 ( .A0(n10481), .A1(n10508), .S(n3403), .Z(N5502) );
  CMXI2X1 U20410 ( .A0(n10488), .A1(n10482), .S(n4118), .Z(n10495) );
  CMX2X1 U20411 ( .A0(n10483), .A1(n10495), .S(n3776), .Z(n10511) );
  CMXI2X1 U20412 ( .A0(n10484), .A1(n10511), .S(n3402), .Z(N5503) );
  CMXI2X1 U20413 ( .A0(n10491), .A1(n10485), .S(n4117), .Z(n10501) );
  CMX2X1 U20414 ( .A0(n10486), .A1(n10501), .S(n3777), .Z(n10514) );
  CMXI2X1 U20415 ( .A0(n10487), .A1(n10514), .S(n3402), .Z(N5504) );
  CMXI2X1 U20416 ( .A0(n10494), .A1(n10488), .S(n4117), .Z(n10504) );
  CMX2X1 U20417 ( .A0(n10489), .A1(n10504), .S(n3790), .Z(n10517) );
  CMXI2X1 U20418 ( .A0(n10490), .A1(n10517), .S(n3402), .Z(N5505) );
  CMXI2X1 U20419 ( .A0(n10500), .A1(n10491), .S(n4117), .Z(n10507) );
  CMX2X1 U20420 ( .A0(n10492), .A1(n10507), .S(n3791), .Z(n10520) );
  CMXI2X1 U20421 ( .A0(n10493), .A1(n10520), .S(n3402), .Z(N5506) );
  CMXI2X1 U20422 ( .A0(n10503), .A1(n10494), .S(n4117), .Z(n10510) );
  CMX2X1 U20423 ( .A0(n10495), .A1(n10510), .S(n3776), .Z(n10523) );
  CMXI2X1 U20424 ( .A0(n10496), .A1(n10523), .S(n3402), .Z(N5507) );
  CMX2X1 U20425 ( .A0(N8231), .A1(N8230), .S(n4256), .Z(n10563) );
  CMXI2X1 U20426 ( .A0(n10563), .A1(n10497), .S(n4117), .Z(n10630) );
  CMX2X1 U20427 ( .A0(n10498), .A1(n10630), .S(n3777), .Z(n10770) );
  CMXI2X1 U20428 ( .A0(n10499), .A1(n10770), .S(n3402), .Z(N5192) );
  CMXI2X1 U20429 ( .A0(n10506), .A1(n10500), .S(n4117), .Z(n10513) );
  CMX2X1 U20430 ( .A0(n10501), .A1(n10513), .S(n3806), .Z(n10526) );
  CMXI2X1 U20431 ( .A0(n10502), .A1(n10526), .S(n3402), .Z(N5508) );
  CMXI2X1 U20432 ( .A0(n10509), .A1(n10503), .S(n4117), .Z(n10516) );
  CMX2X1 U20433 ( .A0(n10504), .A1(n10516), .S(n3791), .Z(n10529) );
  CMXI2X1 U20434 ( .A0(n10505), .A1(n10529), .S(n3301), .Z(N5509) );
  CMXI2X1 U20435 ( .A0(n10512), .A1(n10506), .S(n4117), .Z(n10519) );
  CMX2X1 U20436 ( .A0(n10507), .A1(n10519), .S(n3812), .Z(n10535) );
  CMXI2X1 U20437 ( .A0(n10508), .A1(n10535), .S(n3300), .Z(N5510) );
  CMXI2X1 U20438 ( .A0(n10515), .A1(n10509), .S(n4117), .Z(n10522) );
  CMX2X1 U20439 ( .A0(n10510), .A1(n10522), .S(n3776), .Z(n10538) );
  CMXI2X1 U20440 ( .A0(n10511), .A1(n10538), .S(n3300), .Z(N5511) );
  CMXI2X1 U20441 ( .A0(n10518), .A1(n10512), .S(n4117), .Z(n10525) );
  CMX2X1 U20442 ( .A0(n10513), .A1(n10525), .S(n3772), .Z(n10541) );
  CMXI2X1 U20443 ( .A0(n10514), .A1(n10541), .S(n3300), .Z(N5512) );
  CMXI2X1 U20444 ( .A0(n10521), .A1(n10515), .S(n4117), .Z(n10528) );
  CMX2X1 U20445 ( .A0(n10516), .A1(n10528), .S(n3773), .Z(n10544) );
  CMXI2X1 U20446 ( .A0(n10517), .A1(n10544), .S(n3300), .Z(N5513) );
  CMXI2X1 U20447 ( .A0(n10524), .A1(n10518), .S(n4117), .Z(n10534) );
  CMX2X1 U20448 ( .A0(n10519), .A1(n10534), .S(n3774), .Z(n10547) );
  CMXI2X1 U20449 ( .A0(n10520), .A1(n10547), .S(n3300), .Z(N5514) );
  CMXI2X1 U20450 ( .A0(n10527), .A1(n10521), .S(n4117), .Z(n10537) );
  CMX2X1 U20451 ( .A0(n10522), .A1(n10537), .S(n3775), .Z(n10550) );
  CMXI2X1 U20452 ( .A0(n10523), .A1(n10550), .S(n3300), .Z(N5515) );
  CMXI2X1 U20453 ( .A0(n10533), .A1(n10524), .S(n4117), .Z(n10540) );
  CMX2X1 U20454 ( .A0(n10525), .A1(n10540), .S(n3776), .Z(n10553) );
  CMXI2X1 U20455 ( .A0(n10526), .A1(n10553), .S(n3300), .Z(N5516) );
  CMXI2X1 U20456 ( .A0(n10536), .A1(n10527), .S(n4117), .Z(n10543) );
  CMX2X1 U20457 ( .A0(n10528), .A1(n10543), .S(n3777), .Z(n10556) );
  CMXI2X1 U20458 ( .A0(n10529), .A1(n10556), .S(n3300), .Z(N5517) );
  CMX2X1 U20459 ( .A0(N8230), .A1(N8229), .S(n4260), .Z(n10596) );
  CMXI2X1 U20460 ( .A0(n10596), .A1(n10530), .S(n4117), .Z(n10663) );
  CMX2X1 U20461 ( .A0(n10531), .A1(n10663), .S(n3790), .Z(n10803) );
  CMXI2X1 U20462 ( .A0(n10532), .A1(n10803), .S(n3300), .Z(N5193) );
  CMXI2X1 U20463 ( .A0(n10539), .A1(n10533), .S(n4116), .Z(n10546) );
  CMX2X1 U20464 ( .A0(n10534), .A1(n10546), .S(n3791), .Z(n10559) );
  CMXI2X1 U20465 ( .A0(n10535), .A1(n10559), .S(n3300), .Z(N5518) );
  CMXI2X1 U20466 ( .A0(n10542), .A1(n10536), .S(n4116), .Z(n10549) );
  CMX2X1 U20467 ( .A0(n10537), .A1(n10549), .S(n3792), .Z(n10562) );
  CMXI2X1 U20468 ( .A0(n10538), .A1(n10562), .S(n3412), .Z(N5519) );
  CMXI2X1 U20469 ( .A0(n10545), .A1(n10539), .S(n4116), .Z(n10552) );
  CMX2X1 U20470 ( .A0(n10540), .A1(n10552), .S(n3793), .Z(n10568) );
  CMXI2X1 U20471 ( .A0(n10541), .A1(n10568), .S(n3306), .Z(N5520) );
  CMXI2X1 U20472 ( .A0(n10548), .A1(n10542), .S(n4116), .Z(n10555) );
  CMX2X1 U20473 ( .A0(n10543), .A1(n10555), .S(n3794), .Z(n10571) );
  CMXI2X1 U20474 ( .A0(n10544), .A1(n10571), .S(n3332), .Z(N5521) );
  CMXI2X1 U20475 ( .A0(n10551), .A1(n10545), .S(n4116), .Z(n10558) );
  CMX2X1 U20476 ( .A0(n10546), .A1(n10558), .S(n3795), .Z(n10574) );
  CMXI2X1 U20477 ( .A0(n10547), .A1(n10574), .S(n3332), .Z(N5522) );
  CMXI2X1 U20478 ( .A0(n10554), .A1(n10548), .S(n4116), .Z(n10561) );
  CMX2X1 U20479 ( .A0(n10549), .A1(n10561), .S(n3796), .Z(n10577) );
  CMXI2X1 U20480 ( .A0(n10550), .A1(n10577), .S(n3332), .Z(N5523) );
  CMXI2X1 U20481 ( .A0(n10557), .A1(n10551), .S(n4116), .Z(n10567) );
  CMX2X1 U20482 ( .A0(n10552), .A1(n10567), .S(n3797), .Z(n10580) );
  CMXI2X1 U20483 ( .A0(n10553), .A1(n10580), .S(n3332), .Z(N5524) );
  CMXI2X1 U20484 ( .A0(n10560), .A1(n10554), .S(n4116), .Z(n10570) );
  CMX2X1 U20485 ( .A0(n10555), .A1(n10570), .S(n3805), .Z(n10583) );
  CMXI2X1 U20486 ( .A0(n10556), .A1(n10583), .S(n3332), .Z(N5525) );
  CMXI2X1 U20487 ( .A0(n10566), .A1(n10557), .S(n4116), .Z(n10573) );
  CMX2X1 U20488 ( .A0(n10558), .A1(n10573), .S(n3806), .Z(n10586) );
  CMXI2X1 U20489 ( .A0(n10559), .A1(n10586), .S(n3511), .Z(N5526) );
  CMXI2X1 U20490 ( .A0(n10569), .A1(n10560), .S(n4116), .Z(n10576) );
  CMX2X1 U20491 ( .A0(n10561), .A1(n10576), .S(n3806), .Z(n10589) );
  CMXI2X1 U20492 ( .A0(n10562), .A1(n10589), .S(n3511), .Z(N5527) );
  CMX2X1 U20493 ( .A0(N8229), .A1(N8228), .S(n4259), .Z(n10629) );
  CMXI2X1 U20494 ( .A0(n10629), .A1(n10563), .S(n4116), .Z(n10703) );
  CMX2X1 U20495 ( .A0(n10564), .A1(n10703), .S(n3807), .Z(n10836) );
  CMXI2X1 U20496 ( .A0(n10565), .A1(n10836), .S(n3511), .Z(N5194) );
  CMX2X1 U20497 ( .A0(N7895), .A1(N7894), .S(n4259), .Z(n10572) );
  CMXI2X1 U20498 ( .A0(n10572), .A1(n10566), .S(n4116), .Z(n10579) );
  CMX2X1 U20499 ( .A0(n10567), .A1(n10579), .S(n4317), .Z(n10592) );
  CMXI2X1 U20500 ( .A0(n10568), .A1(n10592), .S(n3511), .Z(N5528) );
  CMX2X1 U20501 ( .A0(N7894), .A1(N7893), .S(n4259), .Z(n10575) );
  CMXI2X1 U20502 ( .A0(n10575), .A1(n10569), .S(n4116), .Z(n10582) );
  CMX2X1 U20503 ( .A0(n10570), .A1(n10582), .S(n3771), .Z(n10595) );
  CMXI2X1 U20504 ( .A0(n10571), .A1(n10595), .S(n3510), .Z(N5529) );
  CMX2X1 U20505 ( .A0(N7893), .A1(N7892), .S(n4259), .Z(n10578) );
  CMXI2X1 U20506 ( .A0(n10578), .A1(n10572), .S(n4116), .Z(n10585) );
  CMX2X1 U20507 ( .A0(n10573), .A1(n10585), .S(n3772), .Z(n10601) );
  CMXI2X1 U20508 ( .A0(n10574), .A1(n10601), .S(n3510), .Z(N5530) );
  CMX2X1 U20509 ( .A0(N7892), .A1(N7891), .S(n4259), .Z(n10581) );
  CMXI2X1 U20510 ( .A0(n10581), .A1(n10575), .S(n4116), .Z(n10588) );
  CMX2X1 U20511 ( .A0(n10576), .A1(n10588), .S(n3773), .Z(n10604) );
  CMXI2X1 U20512 ( .A0(n10577), .A1(n10604), .S(n3510), .Z(N5531) );
  CMX2X1 U20513 ( .A0(N7891), .A1(N7890), .S(n4259), .Z(n10584) );
  CMXI2X1 U20514 ( .A0(n10584), .A1(n10578), .S(n4116), .Z(n10591) );
  CMX2X1 U20515 ( .A0(n10579), .A1(n10591), .S(n3774), .Z(n10607) );
  CMXI2X1 U20516 ( .A0(n10580), .A1(n10607), .S(n3510), .Z(N5532) );
  CMX2X1 U20517 ( .A0(N7890), .A1(N7889), .S(n4258), .Z(n10587) );
  CMXI2X1 U20518 ( .A0(n10587), .A1(n10581), .S(n4115), .Z(n10594) );
  CMX2X1 U20519 ( .A0(n10582), .A1(n10594), .S(n3777), .Z(n10610) );
  CMXI2X1 U20520 ( .A0(n10583), .A1(n10610), .S(n3510), .Z(N5533) );
  CMXI2X1 U20521 ( .A0(n10590), .A1(n10584), .S(n4115), .Z(n10600) );
  CMX2X1 U20522 ( .A0(n10585), .A1(n10600), .S(n3807), .Z(n10613) );
  CMXI2X1 U20523 ( .A0(n10586), .A1(n10613), .S(n3510), .Z(N5534) );
  CMXI2X1 U20524 ( .A0(n10593), .A1(n10587), .S(n4115), .Z(n10603) );
  CMX2X1 U20525 ( .A0(n10588), .A1(n10603), .S(n3808), .Z(n10616) );
  CMXI2X1 U20526 ( .A0(n10589), .A1(n10616), .S(n3510), .Z(N5535) );
  CMX2X1 U20527 ( .A0(N7887), .A1(N7886), .S(n4258), .Z(n10599) );
  CMXI2X1 U20528 ( .A0(n10599), .A1(n10590), .S(n4115), .Z(n10606) );
  CMX2X1 U20529 ( .A0(n10591), .A1(n10606), .S(n3809), .Z(n10619) );
  CMXI2X1 U20530 ( .A0(n10592), .A1(n10619), .S(n3510), .Z(N5536) );
  CMX2X1 U20531 ( .A0(N7886), .A1(N7885), .S(n4258), .Z(n10602) );
  CMXI2X1 U20532 ( .A0(n10602), .A1(n10593), .S(n4115), .Z(n10609) );
  CMX2X1 U20533 ( .A0(n10594), .A1(n10609), .S(n3810), .Z(n10622) );
  CMXI2X1 U20534 ( .A0(n10595), .A1(n10622), .S(n3510), .Z(N5537) );
  CMX2X1 U20535 ( .A0(N8228), .A1(N8227), .S(n4258), .Z(n10662) );
  CMXI2X1 U20536 ( .A0(n10662), .A1(n10596), .S(n4115), .Z(n10736) );
  CMX2X1 U20537 ( .A0(n10597), .A1(n10736), .S(n3811), .Z(n10869) );
  CMXI2X1 U20538 ( .A0(n10598), .A1(n10869), .S(n3510), .Z(N5195) );
  CMXI2X1 U20539 ( .A0(n10605), .A1(n10599), .S(n4115), .Z(n10612) );
  CMX2X1 U20540 ( .A0(n10600), .A1(n10612), .S(n3812), .Z(n10625) );
  CMXI2X1 U20541 ( .A0(n10601), .A1(n10625), .S(n3510), .Z(N5538) );
  CMXI2X1 U20542 ( .A0(n10608), .A1(n10602), .S(n4115), .Z(n10615) );
  CMX2X1 U20543 ( .A0(n10603), .A1(n10615), .S(n4327), .Z(n10628) );
  CMXI2X1 U20544 ( .A0(n10604), .A1(n10628), .S(n3509), .Z(N5539) );
  CMX2X1 U20545 ( .A0(N7883), .A1(N7882), .S(n4258), .Z(n10611) );
  CMXI2X1 U20546 ( .A0(n10611), .A1(n10605), .S(n4115), .Z(n10618) );
  CMX2X1 U20547 ( .A0(n10606), .A1(n10618), .S(n3771), .Z(n10634) );
  CMXI2X1 U20548 ( .A0(n10607), .A1(n10634), .S(n3509), .Z(N5540) );
  CMX2X1 U20549 ( .A0(N7882), .A1(N7881), .S(n4258), .Z(n10614) );
  CMXI2X1 U20550 ( .A0(n10614), .A1(n10608), .S(n4115), .Z(n10621) );
  CMX2X1 U20551 ( .A0(n10609), .A1(n10621), .S(n3772), .Z(n10637) );
  CMXI2X1 U20552 ( .A0(n10610), .A1(n10637), .S(n3509), .Z(N5541) );
  CMXI2X1 U20553 ( .A0(n10617), .A1(n10611), .S(n4115), .Z(n10624) );
  CMX2X1 U20554 ( .A0(n10612), .A1(n10624), .S(n3773), .Z(n10640) );
  CMXI2X1 U20555 ( .A0(n10613), .A1(n10640), .S(n3512), .Z(N5542) );
  CMXI2X1 U20556 ( .A0(n10620), .A1(n10614), .S(n4115), .Z(n10627) );
  CMX2X1 U20557 ( .A0(n10615), .A1(n10627), .S(n3774), .Z(n10643) );
  CMXI2X1 U20558 ( .A0(n10616), .A1(n10643), .S(n3512), .Z(N5543) );
  CMXI2X1 U20559 ( .A0(n10623), .A1(n10617), .S(n4115), .Z(n10633) );
  CMX2X1 U20560 ( .A0(n10618), .A1(n10633), .S(n3775), .Z(n10646) );
  CMXI2X1 U20561 ( .A0(n10619), .A1(n10646), .S(n3512), .Z(N5544) );
  CMXI2X1 U20562 ( .A0(n10626), .A1(n10620), .S(n4115), .Z(n10636) );
  CMX2X1 U20563 ( .A0(n10621), .A1(n10636), .S(n3776), .Z(n10649) );
  CMXI2X1 U20564 ( .A0(n10622), .A1(n10649), .S(n3512), .Z(N5545) );
  CMXI2X1 U20565 ( .A0(n10632), .A1(n10623), .S(n4115), .Z(n10639) );
  CMX2X1 U20566 ( .A0(n10624), .A1(n10639), .S(n3777), .Z(n10652) );
  CMXI2X1 U20567 ( .A0(n10625), .A1(n10652), .S(n3512), .Z(N5546) );
  CMXI2X1 U20568 ( .A0(n10635), .A1(n10626), .S(n4115), .Z(n10642) );
  CMX2X1 U20569 ( .A0(n10627), .A1(n10642), .S(n3790), .Z(n10655) );
  CMXI2X1 U20570 ( .A0(n10628), .A1(n10655), .S(n3512), .Z(N5547) );
  CMX2X1 U20571 ( .A0(N8227), .A1(N8226), .S(n4257), .Z(n10702) );
  CMXI2X1 U20572 ( .A0(n10702), .A1(n10629), .S(n4114), .Z(n10769) );
  CMX2X1 U20573 ( .A0(n10630), .A1(n10769), .S(n3791), .Z(n10902) );
  CMXI2X1 U20574 ( .A0(n10631), .A1(n10902), .S(n3512), .Z(N5196) );
  CMX2X1 U20575 ( .A0(N7875), .A1(N7874), .S(n4257), .Z(n10638) );
  CMXI2X1 U20576 ( .A0(n10638), .A1(n10632), .S(n4114), .Z(n10645) );
  CMX2X1 U20577 ( .A0(n10633), .A1(n10645), .S(n3807), .Z(n10658) );
  CMXI2X1 U20578 ( .A0(n10634), .A1(n10658), .S(n3512), .Z(N5548) );
  CMX2X1 U20579 ( .A0(N7874), .A1(N7873), .S(n4257), .Z(n10641) );
  CMXI2X1 U20580 ( .A0(n10641), .A1(n10635), .S(n4114), .Z(n10648) );
  CMX2X1 U20581 ( .A0(n10636), .A1(n10648), .S(n3808), .Z(n10661) );
  CMXI2X1 U20582 ( .A0(n10637), .A1(n10661), .S(n3512), .Z(N5549) );
  CMX2X1 U20583 ( .A0(N7873), .A1(N7872), .S(n4257), .Z(n10644) );
  CMXI2X1 U20584 ( .A0(n10644), .A1(n10638), .S(n4114), .Z(n10651) );
  CMX2X1 U20585 ( .A0(n10639), .A1(n10651), .S(n3775), .Z(n10674) );
  CMXI2X1 U20586 ( .A0(n10640), .A1(n10674), .S(n3512), .Z(N5550) );
  CMX2X1 U20587 ( .A0(N7872), .A1(N7871), .S(n4257), .Z(n10647) );
  CMXI2X1 U20588 ( .A0(n10647), .A1(n10641), .S(n4114), .Z(n10654) );
  CMX2X1 U20589 ( .A0(n10642), .A1(n10654), .S(n3776), .Z(n10677) );
  CMXI2X1 U20590 ( .A0(n10643), .A1(n10677), .S(n3512), .Z(N5551) );
  CMX2X1 U20591 ( .A0(N7871), .A1(N7870), .S(n4257), .Z(n10650) );
  CMXI2X1 U20592 ( .A0(n10650), .A1(n10644), .S(n4114), .Z(n10657) );
  CMX2X1 U20593 ( .A0(n10645), .A1(n10657), .S(n3777), .Z(n10680) );
  CMXI2X1 U20594 ( .A0(n10646), .A1(n10680), .S(n3511), .Z(N5552) );
  CMX2X1 U20595 ( .A0(N7870), .A1(N7869), .S(n4256), .Z(n10653) );
  CMXI2X1 U20596 ( .A0(n10653), .A1(n10647), .S(n4114), .Z(n10660) );
  CMX2X1 U20597 ( .A0(n10648), .A1(n10660), .S(n3790), .Z(n10683) );
  CMXI2X1 U20598 ( .A0(n10649), .A1(n10683), .S(n3511), .Z(N5553) );
  CMX2X1 U20599 ( .A0(N7869), .A1(N7868), .S(n4256), .Z(n10656) );
  CMXI2X1 U20600 ( .A0(n10656), .A1(n10650), .S(n4114), .Z(n10673) );
  CMX2X1 U20601 ( .A0(n10651), .A1(n10673), .S(n3791), .Z(n10686) );
  CMXI2X1 U20602 ( .A0(n10652), .A1(n10686), .S(n3511), .Z(N5554) );
  CMX2X1 U20603 ( .A0(N7868), .A1(N7867), .S(n4256), .Z(n10659) );
  CMXI2X1 U20604 ( .A0(n10659), .A1(n10653), .S(n4114), .Z(n10676) );
  CMX2X1 U20605 ( .A0(n10654), .A1(n10676), .S(n3790), .Z(n10689) );
  CMXI2X1 U20606 ( .A0(n10655), .A1(n10689), .S(n3511), .Z(N5555) );
  CMXI2X1 U20607 ( .A0(n10672), .A1(n10656), .S(n4114), .Z(n10679) );
  CMX2X1 U20608 ( .A0(n10657), .A1(n10679), .S(n3792), .Z(n10692) );
  CMXI2X1 U20609 ( .A0(n10658), .A1(n10692), .S(n3511), .Z(N5556) );
  CMXI2X1 U20610 ( .A0(n10675), .A1(n10659), .S(n4114), .Z(n10682) );
  CMX2X1 U20611 ( .A0(n10660), .A1(n10682), .S(n3775), .Z(n10695) );
  CMXI2X1 U20612 ( .A0(n10661), .A1(n10695), .S(n3511), .Z(N5557) );
  CMX2X1 U20613 ( .A0(N8226), .A1(N8225), .S(n4256), .Z(n10735) );
  CMXI2X1 U20614 ( .A0(n10735), .A1(n10662), .S(n4114), .Z(n10802) );
  CMX2X1 U20615 ( .A0(n10663), .A1(n10802), .S(n3776), .Z(n10935) );
  CMXI2X1 U20616 ( .A0(n10664), .A1(n10935), .S(n3511), .Z(N5197) );
  CMXI2X1 U20617 ( .A0(n10666), .A1(n10665), .S(n4114), .Z(n12005) );
  CMXI2X1 U20618 ( .A0(n10668), .A1(n10667), .S(n4114), .Z(n10669) );
  CMXI2X1 U20619 ( .A0(n10671), .A1(n10670), .S(n3514), .Z(N5161) );
  CMXI2X1 U20620 ( .A0(n10678), .A1(n10672), .S(n4114), .Z(n10685) );
  CMX2X1 U20621 ( .A0(n10673), .A1(n10685), .S(n3777), .Z(n10698) );
  CMXI2X1 U20622 ( .A0(n10674), .A1(n10698), .S(n3514), .Z(N5558) );
  CMXI2X1 U20623 ( .A0(n10681), .A1(n10675), .S(n4114), .Z(n10688) );
  CMX2X1 U20624 ( .A0(n10676), .A1(n10688), .S(n3790), .Z(n10701) );
  CMXI2X1 U20625 ( .A0(n10677), .A1(n10701), .S(n3514), .Z(N5559) );
  CMXI2X1 U20626 ( .A0(n10684), .A1(n10678), .S(n4113), .Z(n10691) );
  CMX2X1 U20627 ( .A0(n10679), .A1(n10691), .S(n3791), .Z(n10707) );
  CMXI2X1 U20628 ( .A0(n10680), .A1(n10707), .S(n3514), .Z(N5560) );
  CMXI2X1 U20629 ( .A0(n10687), .A1(n10681), .S(n4113), .Z(n10694) );
  CMX2X1 U20630 ( .A0(n10682), .A1(n10694), .S(n3771), .Z(n10710) );
  CMXI2X1 U20631 ( .A0(n10683), .A1(n10710), .S(n3514), .Z(N5561) );
  CMXI2X1 U20632 ( .A0(n10690), .A1(n10684), .S(n4113), .Z(n10697) );
  CMX2X1 U20633 ( .A0(n10685), .A1(n10697), .S(n3807), .Z(n10713) );
  CMXI2X1 U20634 ( .A0(n10686), .A1(n10713), .S(n3514), .Z(N5562) );
  CMXI2X1 U20635 ( .A0(n10693), .A1(n10687), .S(n4113), .Z(n10700) );
  CMX2X1 U20636 ( .A0(n10688), .A1(n10700), .S(n3792), .Z(n10716) );
  CMXI2X1 U20637 ( .A0(n10689), .A1(n10716), .S(n3514), .Z(N5563) );
  CMXI2X1 U20638 ( .A0(n10696), .A1(n10690), .S(n4113), .Z(n10706) );
  CMX2X1 U20639 ( .A0(n10691), .A1(n10706), .S(n3793), .Z(n10719) );
  CMXI2X1 U20640 ( .A0(n10692), .A1(n10719), .S(n3513), .Z(N5564) );
  CMXI2X1 U20641 ( .A0(n10699), .A1(n10693), .S(n4113), .Z(n10709) );
  CMX2X1 U20642 ( .A0(n10694), .A1(n10709), .S(n3794), .Z(n10722) );
  CMXI2X1 U20643 ( .A0(n10695), .A1(n10722), .S(n3513), .Z(N5565) );
  CMXI2X1 U20644 ( .A0(n10705), .A1(n10696), .S(n4113), .Z(n10712) );
  CMX2X1 U20645 ( .A0(n10697), .A1(n10712), .S(n3795), .Z(n10725) );
  CMXI2X1 U20646 ( .A0(n10698), .A1(n10725), .S(n3513), .Z(N5566) );
  CMXI2X1 U20647 ( .A0(n10708), .A1(n10699), .S(n4113), .Z(n10715) );
  CMX2X1 U20648 ( .A0(n10700), .A1(n10715), .S(n3796), .Z(n10728) );
  CMXI2X1 U20649 ( .A0(n10701), .A1(n10728), .S(n3513), .Z(N5567) );
  CMX2X1 U20650 ( .A0(N8225), .A1(N8224), .S(n4248), .Z(n10768) );
  CMXI2X1 U20651 ( .A0(n10768), .A1(n10702), .S(n4113), .Z(n10835) );
  CMX2X1 U20652 ( .A0(n10703), .A1(n10835), .S(n3807), .Z(n10968) );
  CMXI2X1 U20653 ( .A0(n10704), .A1(n10968), .S(n3513), .Z(N5198) );
  CMXI2X1 U20654 ( .A0(n10711), .A1(n10705), .S(n4113), .Z(n10718) );
  CMX2X1 U20655 ( .A0(n10706), .A1(n10718), .S(n3792), .Z(n10731) );
  CMXI2X1 U20656 ( .A0(n10707), .A1(n10731), .S(n3513), .Z(N5568) );
  CMXI2X1 U20657 ( .A0(n10714), .A1(n10708), .S(n4113), .Z(n10721) );
  CMX2X1 U20658 ( .A0(n10709), .A1(n10721), .S(n3793), .Z(n10734) );
  CMXI2X1 U20659 ( .A0(n10710), .A1(n10734), .S(n3513), .Z(N5569) );
  CMXI2X1 U20660 ( .A0(n10717), .A1(n10711), .S(n4113), .Z(n10724) );
  CMX2X1 U20661 ( .A0(n10712), .A1(n10724), .S(n3794), .Z(n10740) );
  CMXI2X1 U20662 ( .A0(n10713), .A1(n10740), .S(n3513), .Z(N5570) );
  CMXI2X1 U20663 ( .A0(n10720), .A1(n10714), .S(n4113), .Z(n10727) );
  CMX2X1 U20664 ( .A0(n10715), .A1(n10727), .S(n3795), .Z(n10743) );
  CMXI2X1 U20665 ( .A0(n10716), .A1(n10743), .S(n3513), .Z(N5571) );
  CMXI2X1 U20666 ( .A0(n10723), .A1(n10717), .S(n4113), .Z(n10730) );
  CMX2X1 U20667 ( .A0(n10718), .A1(n10730), .S(n3796), .Z(n10746) );
  CMXI2X1 U20668 ( .A0(n10719), .A1(n10746), .S(n3513), .Z(N5572) );
  CMXI2X1 U20669 ( .A0(n10726), .A1(n10720), .S(n4113), .Z(n10733) );
  CMX2X1 U20670 ( .A0(n10721), .A1(n10733), .S(n3797), .Z(n10749) );
  CMXI2X1 U20671 ( .A0(n10722), .A1(n10749), .S(n3513), .Z(N5573) );
  CMXI2X1 U20672 ( .A0(n10729), .A1(n10723), .S(n4113), .Z(n10739) );
  CMX2X1 U20673 ( .A0(n10724), .A1(n10739), .S(n3805), .Z(n10752) );
  CMXI2X1 U20674 ( .A0(n10725), .A1(n10752), .S(n3412), .Z(N5574) );
  CMXI2X1 U20675 ( .A0(n10732), .A1(n10726), .S(n4112), .Z(n10742) );
  CMX2X1 U20676 ( .A0(n10727), .A1(n10742), .S(n3806), .Z(n10755) );
  CMXI2X1 U20677 ( .A0(n10728), .A1(n10755), .S(n3412), .Z(N5575) );
  CMXI2X1 U20678 ( .A0(n10738), .A1(n10729), .S(n4112), .Z(n10745) );
  CMX2X1 U20679 ( .A0(n10730), .A1(n10745), .S(n3807), .Z(n10758) );
  CMXI2X1 U20680 ( .A0(n10731), .A1(n10758), .S(n3412), .Z(N5576) );
  CMXI2X1 U20681 ( .A0(n10741), .A1(n10732), .S(n4112), .Z(n10748) );
  CMX2X1 U20682 ( .A0(n10733), .A1(n10748), .S(n3809), .Z(n10761) );
  CMXI2X1 U20683 ( .A0(n10734), .A1(n10761), .S(n3420), .Z(N5577) );
  CMX2X1 U20684 ( .A0(N8224), .A1(N8223), .S(n4228), .Z(n10801) );
  CMXI2X1 U20685 ( .A0(n10801), .A1(n10735), .S(n4112), .Z(n10868) );
  CMX2X1 U20686 ( .A0(n10736), .A1(n10868), .S(n3810), .Z(n11001) );
  CMXI2X1 U20687 ( .A0(n10737), .A1(n11001), .S(n3429), .Z(N5199) );
  CMXI2X1 U20688 ( .A0(n10744), .A1(n10738), .S(n4112), .Z(n10751) );
  CMX2X1 U20689 ( .A0(n10739), .A1(n10751), .S(n3811), .Z(n10764) );
  CMXI2X1 U20690 ( .A0(n10740), .A1(n10764), .S(n3515), .Z(N5578) );
  CMXI2X1 U20691 ( .A0(n10747), .A1(n10741), .S(n4112), .Z(n10754) );
  CMX2X1 U20692 ( .A0(n10742), .A1(n10754), .S(n3771), .Z(n10767) );
  CMXI2X1 U20693 ( .A0(n10743), .A1(n10767), .S(n3515), .Z(N5579) );
  CMXI2X1 U20694 ( .A0(n10750), .A1(n10744), .S(n4112), .Z(n10757) );
  CMX2X1 U20695 ( .A0(n10745), .A1(n10757), .S(n3807), .Z(n10773) );
  CMXI2X1 U20696 ( .A0(n10746), .A1(n10773), .S(n3515), .Z(N5580) );
  CMXI2X1 U20697 ( .A0(n10753), .A1(n10747), .S(n4112), .Z(n10760) );
  CMX2X1 U20698 ( .A0(n10748), .A1(n10760), .S(n3808), .Z(n10776) );
  CMXI2X1 U20699 ( .A0(n10749), .A1(n10776), .S(n3515), .Z(N5581) );
  CMXI2X1 U20700 ( .A0(n10756), .A1(n10750), .S(n4112), .Z(n10763) );
  CMX2X1 U20701 ( .A0(n10751), .A1(n10763), .S(n3809), .Z(n10779) );
  CMXI2X1 U20702 ( .A0(n10752), .A1(n10779), .S(n3515), .Z(N5582) );
  CMXI2X1 U20703 ( .A0(n10759), .A1(n10753), .S(n4112), .Z(n10766) );
  CMX2X1 U20704 ( .A0(n10754), .A1(n10766), .S(n3810), .Z(n10782) );
  CMXI2X1 U20705 ( .A0(n10755), .A1(n10782), .S(n3515), .Z(N5583) );
  CMXI2X1 U20706 ( .A0(n10762), .A1(n10756), .S(n4112), .Z(n10772) );
  CMX2X1 U20707 ( .A0(n10757), .A1(n10772), .S(n3811), .Z(n10785) );
  CMXI2X1 U20708 ( .A0(n10758), .A1(n10785), .S(n3515), .Z(N5584) );
  CMXI2X1 U20709 ( .A0(n10765), .A1(n10759), .S(n4112), .Z(n10775) );
  CMX2X1 U20710 ( .A0(n10760), .A1(n10775), .S(n3812), .Z(n10788) );
  CMXI2X1 U20711 ( .A0(n10761), .A1(n10788), .S(n3515), .Z(N5585) );
  CMXI2X1 U20712 ( .A0(n10771), .A1(n10762), .S(n4112), .Z(n10778) );
  CMX2X1 U20713 ( .A0(n10763), .A1(n10778), .S(n4333), .Z(n10791) );
  CMXI2X1 U20714 ( .A0(n10764), .A1(n10791), .S(n3515), .Z(N5586) );
  CMXI2X1 U20715 ( .A0(n10774), .A1(n10765), .S(n4112), .Z(n10781) );
  CMX2X1 U20716 ( .A0(n10766), .A1(n10781), .S(n3771), .Z(n10794) );
  CMXI2X1 U20717 ( .A0(n10767), .A1(n10794), .S(n3514), .Z(N5587) );
  CMX2X1 U20718 ( .A0(N8223), .A1(N8222), .S(n4236), .Z(n10834) );
  CMXI2X1 U20719 ( .A0(n10834), .A1(n10768), .S(n4112), .Z(n10901) );
  CMX2X1 U20720 ( .A0(n10769), .A1(n10901), .S(n3772), .Z(n11038) );
  CMXI2X1 U20721 ( .A0(n10770), .A1(n11038), .S(n3514), .Z(N5200) );
  CMXI2X1 U20722 ( .A0(n10777), .A1(n10771), .S(n4112), .Z(n10784) );
  CMX2X1 U20723 ( .A0(n10772), .A1(n10784), .S(n3773), .Z(n10797) );
  CMXI2X1 U20724 ( .A0(n10773), .A1(n10797), .S(n3514), .Z(N5588) );
  CMXI2X1 U20725 ( .A0(n10780), .A1(n10774), .S(n4111), .Z(n10787) );
  CMX2X1 U20726 ( .A0(n10775), .A1(n10787), .S(n3774), .Z(n10800) );
  CMXI2X1 U20727 ( .A0(n10776), .A1(n10800), .S(n3514), .Z(N5589) );
  CMXI2X1 U20728 ( .A0(n10783), .A1(n10777), .S(n4111), .Z(n10790) );
  CMX2X1 U20729 ( .A0(n10778), .A1(n10790), .S(n3775), .Z(n10806) );
  CMXI2X1 U20730 ( .A0(n10779), .A1(n10806), .S(n3413), .Z(N5590) );
  CMXI2X1 U20731 ( .A0(n10786), .A1(n10780), .S(n4111), .Z(n10793) );
  CMX2X1 U20732 ( .A0(n10781), .A1(n10793), .S(n3776), .Z(n10809) );
  CMXI2X1 U20733 ( .A0(n10782), .A1(n10809), .S(n3413), .Z(N5591) );
  CMX2X1 U20734 ( .A0(N7831), .A1(N7830), .S(n4255), .Z(n10789) );
  CMXI2X1 U20735 ( .A0(n10789), .A1(n10783), .S(n4111), .Z(n10796) );
  CMX2X1 U20736 ( .A0(n10784), .A1(n10796), .S(n3777), .Z(n10812) );
  CMXI2X1 U20737 ( .A0(n10785), .A1(n10812), .S(n3413), .Z(N5592) );
  CMX2X1 U20738 ( .A0(N7830), .A1(N7829), .S(n4255), .Z(n10792) );
  CMXI2X1 U20739 ( .A0(n10792), .A1(n10786), .S(n4111), .Z(n10799) );
  CMX2X1 U20740 ( .A0(n10787), .A1(n10799), .S(n3790), .Z(n10815) );
  CMXI2X1 U20741 ( .A0(n10788), .A1(n10815), .S(n3413), .Z(N5593) );
  CMX2X1 U20742 ( .A0(N7829), .A1(N7828), .S(n4255), .Z(n10795) );
  CMXI2X1 U20743 ( .A0(n10795), .A1(n10789), .S(n4111), .Z(n10805) );
  CMX2X1 U20744 ( .A0(n10790), .A1(n10805), .S(n3791), .Z(n10818) );
  CMXI2X1 U20745 ( .A0(n10791), .A1(n10818), .S(n3413), .Z(N5594) );
  CMX2X1 U20746 ( .A0(N7828), .A1(N7827), .S(n4255), .Z(n10798) );
  CMXI2X1 U20747 ( .A0(n10798), .A1(n10792), .S(n4111), .Z(n10808) );
  CMX2X1 U20748 ( .A0(n10793), .A1(n10808), .S(n3794), .Z(n10821) );
  CMXI2X1 U20749 ( .A0(n10794), .A1(n10821), .S(n3413), .Z(N5595) );
  CMXI2X1 U20750 ( .A0(n10804), .A1(n10795), .S(n4111), .Z(n10811) );
  CMX2X1 U20751 ( .A0(n10796), .A1(n10811), .S(n3812), .Z(n10824) );
  CMXI2X1 U20752 ( .A0(n10797), .A1(n10824), .S(n3413), .Z(N5596) );
  CMXI2X1 U20753 ( .A0(n10807), .A1(n10798), .S(n4111), .Z(n10814) );
  CMX2X1 U20754 ( .A0(n10799), .A1(n10814), .S(n4318), .Z(n10827) );
  CMXI2X1 U20755 ( .A0(n10800), .A1(n10827), .S(n3413), .Z(N5597) );
  CMX2X1 U20756 ( .A0(N8222), .A1(N8221), .S(n4255), .Z(n10867) );
  CMXI2X1 U20757 ( .A0(n10867), .A1(n10801), .S(n4111), .Z(n10934) );
  CMX2X1 U20758 ( .A0(n10802), .A1(n10934), .S(n3771), .Z(n11071) );
  CMXI2X1 U20759 ( .A0(n10803), .A1(n11071), .S(n3413), .Z(N5201) );
  CMXI2X1 U20760 ( .A0(n10810), .A1(n10804), .S(n4111), .Z(n10817) );
  CMX2X1 U20761 ( .A0(n10805), .A1(n10817), .S(n3772), .Z(n10830) );
  CMXI2X1 U20762 ( .A0(n10806), .A1(n10830), .S(n3413), .Z(N5598) );
  CMXI2X1 U20763 ( .A0(n10813), .A1(n10807), .S(n4111), .Z(n10820) );
  CMX2X1 U20764 ( .A0(n10808), .A1(n10820), .S(n3773), .Z(n10833) );
  CMXI2X1 U20765 ( .A0(n10809), .A1(n10833), .S(n3412), .Z(N5599) );
  CMX2X1 U20766 ( .A0(N7823), .A1(N7822), .S(n4255), .Z(n10816) );
  CMXI2X1 U20767 ( .A0(n10816), .A1(n10810), .S(n4111), .Z(n10823) );
  CMX2X1 U20768 ( .A0(n10811), .A1(n10823), .S(n3772), .Z(n10839) );
  CMXI2X1 U20769 ( .A0(n10812), .A1(n10839), .S(n3412), .Z(N5600) );
  CMX2X1 U20770 ( .A0(N7822), .A1(N7821), .S(n4255), .Z(n10819) );
  CMXI2X1 U20771 ( .A0(n10819), .A1(n10813), .S(n4111), .Z(n10826) );
  CMX2X1 U20772 ( .A0(n10814), .A1(n10826), .S(n3792), .Z(n10842) );
  CMXI2X1 U20773 ( .A0(n10815), .A1(n10842), .S(n3412), .Z(N5601) );
  CMX2X1 U20774 ( .A0(N7821), .A1(N7820), .S(n4254), .Z(n10822) );
  CMXI2X1 U20775 ( .A0(n10822), .A1(n10816), .S(n4111), .Z(n10829) );
  CMX2X1 U20776 ( .A0(n10817), .A1(n10829), .S(n3793), .Z(n10845) );
  CMXI2X1 U20777 ( .A0(n10818), .A1(n10845), .S(n3412), .Z(N5602) );
  CMX2X1 U20778 ( .A0(N7820), .A1(N7819), .S(n4254), .Z(n10825) );
  CMXI2X1 U20779 ( .A0(n10825), .A1(n10819), .S(n4111), .Z(n10832) );
  CMX2X1 U20780 ( .A0(n10820), .A1(n10832), .S(n3794), .Z(n10848) );
  CMXI2X1 U20781 ( .A0(n10821), .A1(n10848), .S(n3412), .Z(N5603) );
  CMX2X1 U20782 ( .A0(N7819), .A1(N7818), .S(n4254), .Z(n10828) );
  CMXI2X1 U20783 ( .A0(n10828), .A1(n10822), .S(n4110), .Z(n10838) );
  CMX2X1 U20784 ( .A0(n10823), .A1(n10838), .S(n3795), .Z(n10851) );
  CMXI2X1 U20785 ( .A0(n10824), .A1(n10851), .S(n3412), .Z(N5604) );
  CMX2X1 U20786 ( .A0(N7818), .A1(N7817), .S(n4254), .Z(n10831) );
  CMXI2X1 U20787 ( .A0(n10831), .A1(n10825), .S(n4110), .Z(n10841) );
  CMX2X1 U20788 ( .A0(n10826), .A1(n10841), .S(n3796), .Z(n10854) );
  CMXI2X1 U20789 ( .A0(n10827), .A1(n10854), .S(n3412), .Z(N5605) );
  CMXI2X1 U20790 ( .A0(n10837), .A1(n10828), .S(n4110), .Z(n10844) );
  CMX2X1 U20791 ( .A0(n10829), .A1(n10844), .S(n3797), .Z(n10857) );
  CMXI2X1 U20792 ( .A0(n10830), .A1(n10857), .S(n3415), .Z(N5606) );
  CMXI2X1 U20793 ( .A0(n10840), .A1(n10831), .S(n4110), .Z(n10847) );
  CMX2X1 U20794 ( .A0(n10832), .A1(n10847), .S(n3805), .Z(n10860) );
  CMXI2X1 U20795 ( .A0(n10833), .A1(n10860), .S(n3415), .Z(N5607) );
  CMX2X1 U20796 ( .A0(N8221), .A1(N8220), .S(n4254), .Z(n10900) );
  CMXI2X1 U20797 ( .A0(n10900), .A1(n10834), .S(n4110), .Z(n10967) );
  CMX2X1 U20798 ( .A0(n10835), .A1(n10967), .S(n3806), .Z(n11104) );
  CMXI2X1 U20799 ( .A0(n10836), .A1(n11104), .S(n3415), .Z(N5202) );
  CMXI2X1 U20800 ( .A0(n10843), .A1(n10837), .S(n4110), .Z(n10850) );
  CMX2X1 U20801 ( .A0(n10838), .A1(n10850), .S(n3807), .Z(n10863) );
  CMXI2X1 U20802 ( .A0(n10839), .A1(n10863), .S(n3415), .Z(N5608) );
  CMXI2X1 U20803 ( .A0(n10846), .A1(n10840), .S(n4110), .Z(n10853) );
  CMX2X1 U20804 ( .A0(n10841), .A1(n10853), .S(n3808), .Z(n10866) );
  CMXI2X1 U20805 ( .A0(n10842), .A1(n10866), .S(n3415), .Z(N5609) );
  CMX2X1 U20806 ( .A0(N7813), .A1(N7812), .S(n4254), .Z(n10849) );
  CMXI2X1 U20807 ( .A0(n10849), .A1(n10843), .S(n4110), .Z(n10856) );
  CMX2X1 U20808 ( .A0(n10844), .A1(n10856), .S(n3809), .Z(n10872) );
  CMXI2X1 U20809 ( .A0(n10845), .A1(n10872), .S(n3415), .Z(N5610) );
  CMX2X1 U20810 ( .A0(N7812), .A1(N7811), .S(n4254), .Z(n10852) );
  CMXI2X1 U20811 ( .A0(n10852), .A1(n10846), .S(n4110), .Z(n10859) );
  CMX2X1 U20812 ( .A0(n10847), .A1(n10859), .S(n3810), .Z(n10875) );
  CMXI2X1 U20813 ( .A0(n10848), .A1(n10875), .S(n3414), .Z(N5611) );
  CMX2X1 U20814 ( .A0(N7811), .A1(N7810), .S(n4253), .Z(n10855) );
  CMXI2X1 U20815 ( .A0(n10855), .A1(n10849), .S(n4110), .Z(n10862) );
  CMX2X1 U20816 ( .A0(n10850), .A1(n10862), .S(n3811), .Z(n10878) );
  CMXI2X1 U20817 ( .A0(n10851), .A1(n10878), .S(n3414), .Z(N5612) );
  CMX2X1 U20818 ( .A0(N7810), .A1(N7809), .S(n4253), .Z(n10858) );
  CMXI2X1 U20819 ( .A0(n10858), .A1(n10852), .S(n4110), .Z(n10865) );
  CMX2X1 U20820 ( .A0(n10853), .A1(n10865), .S(n3812), .Z(n10881) );
  CMXI2X1 U20821 ( .A0(n10854), .A1(n10881), .S(n3414), .Z(N5613) );
  CMX2X1 U20822 ( .A0(N7809), .A1(N7808), .S(n4253), .Z(n10861) );
  CMXI2X1 U20823 ( .A0(n10861), .A1(n10855), .S(n4110), .Z(n10871) );
  CMX2X1 U20824 ( .A0(n10856), .A1(n10871), .S(n4332), .Z(n10884) );
  CMXI2X1 U20825 ( .A0(n10857), .A1(n10884), .S(n3414), .Z(N5614) );
  CMX2X1 U20826 ( .A0(N7808), .A1(N7807), .S(n4253), .Z(n10864) );
  CMXI2X1 U20827 ( .A0(n10864), .A1(n10858), .S(n4110), .Z(n10874) );
  CMX2X1 U20828 ( .A0(n10859), .A1(n10874), .S(n3771), .Z(n10887) );
  CMXI2X1 U20829 ( .A0(n10860), .A1(n10887), .S(n3414), .Z(N5615) );
  CMX2X1 U20830 ( .A0(N7807), .A1(N7806), .S(n4253), .Z(n10870) );
  CMXI2X1 U20831 ( .A0(n10870), .A1(n10861), .S(n4110), .Z(n10877) );
  CMX2X1 U20832 ( .A0(n10862), .A1(n10877), .S(n3795), .Z(n10890) );
  CMXI2X1 U20833 ( .A0(n10863), .A1(n10890), .S(n3414), .Z(N5616) );
  CMX2X1 U20834 ( .A0(N7806), .A1(N7805), .S(n4253), .Z(n10873) );
  CMXI2X1 U20835 ( .A0(n10873), .A1(n10864), .S(n4110), .Z(n10880) );
  CMX2X1 U20836 ( .A0(n10865), .A1(n10880), .S(n3796), .Z(n10893) );
  CMXI2X1 U20837 ( .A0(n10866), .A1(n10893), .S(n3414), .Z(N5617) );
  CMXI2X1 U20838 ( .A0(n10933), .A1(n10867), .S(n4110), .Z(n11000) );
  CMX2X1 U20839 ( .A0(n10868), .A1(n11000), .S(n3774), .Z(n11137) );
  CMXI2X1 U20840 ( .A0(n10869), .A1(n11137), .S(n3414), .Z(N5203) );
  CMX2X1 U20841 ( .A0(N7805), .A1(N7804), .S(n4253), .Z(n10876) );
  CMXI2X1 U20842 ( .A0(n10876), .A1(n10870), .S(n4109), .Z(n10883) );
  CMX2X1 U20843 ( .A0(n10871), .A1(n10883), .S(n3775), .Z(n10896) );
  CMXI2X1 U20844 ( .A0(n10872), .A1(n10896), .S(n3414), .Z(N5618) );
  CMX2X1 U20845 ( .A0(N7804), .A1(N7803), .S(n4253), .Z(n10879) );
  CMXI2X1 U20846 ( .A0(n10879), .A1(n10873), .S(n4109), .Z(n10886) );
  CMX2X1 U20847 ( .A0(n10874), .A1(n10886), .S(n3776), .Z(n10899) );
  CMXI2X1 U20848 ( .A0(n10875), .A1(n10899), .S(n3414), .Z(N5619) );
  CMXI2X1 U20849 ( .A0(n10882), .A1(n10876), .S(n4109), .Z(n10889) );
  CMX2X1 U20850 ( .A0(n10877), .A1(n10889), .S(n3777), .Z(n10905) );
  CMXI2X1 U20851 ( .A0(n10878), .A1(n10905), .S(n3414), .Z(N5620) );
  CMXI2X1 U20852 ( .A0(n10885), .A1(n10879), .S(n4109), .Z(n10892) );
  CMX2X1 U20853 ( .A0(n10880), .A1(n10892), .S(n3790), .Z(n10908) );
  CMXI2X1 U20854 ( .A0(n10881), .A1(n10908), .S(n3413), .Z(N5621) );
  CMX2X1 U20855 ( .A0(N7801), .A1(N7800), .S(n4229), .Z(n10888) );
  CMXI2X1 U20856 ( .A0(n10888), .A1(n10882), .S(n4109), .Z(n10895) );
  CMX2X1 U20857 ( .A0(n10883), .A1(n10895), .S(n3773), .Z(n10911) );
  CMXI2X1 U20858 ( .A0(n10884), .A1(n10911), .S(n3417), .Z(N5622) );
  CMX2X1 U20859 ( .A0(N7800), .A1(N7799), .S(n4230), .Z(n10891) );
  CMXI2X1 U20860 ( .A0(n10891), .A1(n10885), .S(n4109), .Z(n10898) );
  CMX2X1 U20861 ( .A0(n10886), .A1(n10898), .S(n3772), .Z(n10914) );
  CMXI2X1 U20862 ( .A0(n10887), .A1(n10914), .S(n3417), .Z(N5623) );
  CMXI2X1 U20863 ( .A0(n10894), .A1(n10888), .S(n4109), .Z(n10904) );
  CMX2X1 U20864 ( .A0(n10889), .A1(n10904), .S(n3773), .Z(n10917) );
  CMXI2X1 U20865 ( .A0(n10890), .A1(n10917), .S(n3416), .Z(N5624) );
  CMXI2X1 U20866 ( .A0(n10897), .A1(n10891), .S(n4109), .Z(n10907) );
  CMX2X1 U20867 ( .A0(n10892), .A1(n10907), .S(n3774), .Z(n10920) );
  CMXI2X1 U20868 ( .A0(n10893), .A1(n10920), .S(n3416), .Z(N5625) );
  CMXI2X1 U20869 ( .A0(n10903), .A1(n10894), .S(n4109), .Z(n10910) );
  CMX2X1 U20870 ( .A0(n10895), .A1(n10910), .S(n3775), .Z(n10923) );
  CMXI2X1 U20871 ( .A0(n10896), .A1(n10923), .S(n3416), .Z(N5626) );
  CMXI2X1 U20872 ( .A0(n10906), .A1(n10897), .S(n4109), .Z(n10913) );
  CMX2X1 U20873 ( .A0(n10898), .A1(n10913), .S(n3776), .Z(n10926) );
  CMXI2X1 U20874 ( .A0(n10899), .A1(n10926), .S(n3416), .Z(N5627) );
  CMXI2X1 U20875 ( .A0(n10966), .A1(n10900), .S(n4109), .Z(n11037) );
  CMX2X1 U20876 ( .A0(n10901), .A1(n11037), .S(n3777), .Z(n11170) );
  CMXI2X1 U20877 ( .A0(n10902), .A1(n11170), .S(n3416), .Z(N5204) );
  CMXI2X1 U20878 ( .A0(n10909), .A1(n10903), .S(n4109), .Z(n10916) );
  CMX2X1 U20879 ( .A0(n10904), .A1(n10916), .S(n3790), .Z(n10929) );
  CMXI2X1 U20880 ( .A0(n10905), .A1(n10929), .S(n3416), .Z(N5628) );
  CMXI2X1 U20881 ( .A0(n10912), .A1(n10906), .S(n4109), .Z(n10919) );
  CMX2X1 U20882 ( .A0(n10907), .A1(n10919), .S(n3791), .Z(n10932) );
  CMXI2X1 U20883 ( .A0(n10908), .A1(n10932), .S(n3416), .Z(N5629) );
  CMXI2X1 U20884 ( .A0(n10915), .A1(n10909), .S(n4109), .Z(n10922) );
  CMX2X1 U20885 ( .A0(n10910), .A1(n10922), .S(n3792), .Z(n10938) );
  CMXI2X1 U20886 ( .A0(n10911), .A1(n10938), .S(n3416), .Z(N5630) );
  CMXI2X1 U20887 ( .A0(n10918), .A1(n10912), .S(n4109), .Z(n10925) );
  CMX2X1 U20888 ( .A0(n10913), .A1(n10925), .S(n3793), .Z(n10941) );
  CMXI2X1 U20889 ( .A0(n10914), .A1(n10941), .S(n3416), .Z(N5631) );
  CMXI2X1 U20890 ( .A0(n10921), .A1(n10915), .S(n4109), .Z(n10928) );
  CMX2X1 U20891 ( .A0(n10916), .A1(n10928), .S(n3794), .Z(n10944) );
  CMXI2X1 U20892 ( .A0(n10917), .A1(n10944), .S(n3416), .Z(N5632) );
  CMXI2X1 U20893 ( .A0(n10924), .A1(n10918), .S(n4108), .Z(n10931) );
  CMX2X1 U20894 ( .A0(n10919), .A1(n10931), .S(n3795), .Z(n10947) );
  CMXI2X1 U20895 ( .A0(n10920), .A1(n10947), .S(n3416), .Z(N5633) );
  CMXI2X1 U20896 ( .A0(n10927), .A1(n10921), .S(n4108), .Z(n10937) );
  CMX2X1 U20897 ( .A0(n10922), .A1(n10937), .S(n3796), .Z(n10950) );
  CMXI2X1 U20898 ( .A0(n10923), .A1(n10950), .S(n3415), .Z(N5634) );
  CMXI2X1 U20899 ( .A0(n10930), .A1(n10924), .S(n4108), .Z(n10940) );
  CMX2X1 U20900 ( .A0(n10925), .A1(n10940), .S(n3797), .Z(n10953) );
  CMXI2X1 U20901 ( .A0(n10926), .A1(n10953), .S(n3415), .Z(N5635) );
  CMXI2X1 U20902 ( .A0(n10936), .A1(n10927), .S(n4108), .Z(n10943) );
  CMX2X1 U20903 ( .A0(n10928), .A1(n10943), .S(n3805), .Z(n10956) );
  CMXI2X1 U20904 ( .A0(n10929), .A1(n10956), .S(n3415), .Z(N5636) );
  CMXI2X1 U20905 ( .A0(n10939), .A1(n10930), .S(n4108), .Z(n10946) );
  CMX2X1 U20906 ( .A0(n10931), .A1(n10946), .S(n3806), .Z(n10959) );
  CMXI2X1 U20907 ( .A0(n10932), .A1(n10959), .S(n3415), .Z(N5637) );
  CMXI2X1 U20908 ( .A0(n10999), .A1(n10933), .S(n4108), .Z(n11070) );
  CMX2X1 U20909 ( .A0(n10934), .A1(n11070), .S(n3796), .Z(n11203) );
  CMXI2X1 U20910 ( .A0(n10935), .A1(n11203), .S(n3415), .Z(N5205) );
  CMXI2X1 U20911 ( .A0(n10942), .A1(n10936), .S(n4108), .Z(n10949) );
  CMX2X1 U20912 ( .A0(n10937), .A1(n10949), .S(n3797), .Z(n10962) );
  CMXI2X1 U20913 ( .A0(n10938), .A1(n10962), .S(n3418), .Z(N5638) );
  CMXI2X1 U20914 ( .A0(n10945), .A1(n10939), .S(n4108), .Z(n10952) );
  CMX2X1 U20915 ( .A0(n10940), .A1(n10952), .S(n3791), .Z(n10965) );
  CMXI2X1 U20916 ( .A0(n10941), .A1(n10965), .S(n3418), .Z(N5639) );
  CMXI2X1 U20917 ( .A0(n10948), .A1(n10942), .S(n4108), .Z(n10955) );
  CMX2X1 U20918 ( .A0(n10943), .A1(n10955), .S(n3792), .Z(n10971) );
  CMXI2X1 U20919 ( .A0(n10944), .A1(n10971), .S(n3418), .Z(N5640) );
  CMX2X1 U20920 ( .A0(N7782), .A1(N7781), .S(n4260), .Z(n10951) );
  CMXI2X1 U20921 ( .A0(n10951), .A1(n10945), .S(n4108), .Z(n10958) );
  CMX2X1 U20922 ( .A0(n10946), .A1(n10958), .S(n3793), .Z(n10974) );
  CMXI2X1 U20923 ( .A0(n10947), .A1(n10974), .S(n3418), .Z(N5641) );
  CMXI2X1 U20924 ( .A0(n10954), .A1(n10948), .S(n4108), .Z(n10961) );
  CMX2X1 U20925 ( .A0(n10949), .A1(n10961), .S(n3794), .Z(n10977) );
  CMXI2X1 U20926 ( .A0(n10950), .A1(n10977), .S(n3418), .Z(N5642) );
  CMXI2X1 U20927 ( .A0(n10957), .A1(n10951), .S(n4108), .Z(n10964) );
  CMX2X1 U20928 ( .A0(n10952), .A1(n10964), .S(n3795), .Z(n10980) );
  CMXI2X1 U20929 ( .A0(n10953), .A1(n10980), .S(n3418), .Z(N5643) );
  CMX2X1 U20930 ( .A0(N7779), .A1(N7778), .S(n4252), .Z(n10960) );
  CMXI2X1 U20931 ( .A0(n10960), .A1(n10954), .S(n4108), .Z(n10970) );
  CMX2X1 U20932 ( .A0(n10955), .A1(n10970), .S(n3774), .Z(n10983) );
  CMXI2X1 U20933 ( .A0(n10956), .A1(n10983), .S(n3418), .Z(N5644) );
  CMX2X1 U20934 ( .A0(N7778), .A1(N7777), .S(n4252), .Z(n10963) );
  CMXI2X1 U20935 ( .A0(n10963), .A1(n10957), .S(n4108), .Z(n10973) );
  CMX2X1 U20936 ( .A0(n10958), .A1(n10973), .S(n3807), .Z(n10986) );
  CMXI2X1 U20937 ( .A0(n10959), .A1(n10986), .S(n3418), .Z(N5645) );
  CMX2X1 U20938 ( .A0(N7777), .A1(N7776), .S(n4252), .Z(n10969) );
  CMXI2X1 U20939 ( .A0(n10969), .A1(n10960), .S(n4108), .Z(n10976) );
  CMX2X1 U20940 ( .A0(n10961), .A1(n10976), .S(n3808), .Z(n10989) );
  CMXI2X1 U20941 ( .A0(n10962), .A1(n10989), .S(n3418), .Z(N5646) );
  CMX2X1 U20942 ( .A0(N7776), .A1(N7775), .S(n4252), .Z(n10972) );
  CMXI2X1 U20943 ( .A0(n10972), .A1(n10963), .S(n4108), .Z(n10979) );
  CMX2X1 U20944 ( .A0(n10964), .A1(n10979), .S(n3809), .Z(n10992) );
  CMXI2X1 U20945 ( .A0(n10965), .A1(n10992), .S(n3417), .Z(N5647) );
  CMXI2X1 U20946 ( .A0(n11036), .A1(n10966), .S(n4107), .Z(n11103) );
  CMX2X1 U20947 ( .A0(n10967), .A1(n11103), .S(n3810), .Z(n11236) );
  CMXI2X1 U20948 ( .A0(n10968), .A1(n11236), .S(n3417), .Z(N5206) );
  CMX2X1 U20949 ( .A0(N7775), .A1(N7774), .S(n4252), .Z(n10975) );
  CMXI2X1 U20950 ( .A0(n10975), .A1(n10969), .S(n4107), .Z(n10982) );
  CMX2X1 U20951 ( .A0(n10970), .A1(n10982), .S(n3811), .Z(n10995) );
  CMXI2X1 U20952 ( .A0(n10971), .A1(n10995), .S(n3417), .Z(N5648) );
  CMX2X1 U20953 ( .A0(N7774), .A1(N7773), .S(n4252), .Z(n10978) );
  CMXI2X1 U20954 ( .A0(n10978), .A1(n10972), .S(n4107), .Z(n10985) );
  CMX2X1 U20955 ( .A0(n10973), .A1(n10985), .S(n3812), .Z(n10998) );
  CMXI2X1 U20956 ( .A0(n10974), .A1(n10998), .S(n3417), .Z(N5649) );
  CMX2X1 U20957 ( .A0(N7773), .A1(N7772), .S(n4252), .Z(n10981) );
  CMXI2X1 U20958 ( .A0(n10981), .A1(n10975), .S(n4107), .Z(n10988) );
  CMX2X1 U20959 ( .A0(n10976), .A1(n10988), .S(n4331), .Z(n11008) );
  CMXI2X1 U20960 ( .A0(n10977), .A1(n11008), .S(n3417), .Z(N5650) );
  CMX2X1 U20961 ( .A0(N7772), .A1(N7771), .S(n4252), .Z(n10984) );
  CMXI2X1 U20962 ( .A0(n10984), .A1(n10978), .S(n4107), .Z(n10991) );
  CMX2X1 U20963 ( .A0(n10979), .A1(n10991), .S(n3771), .Z(n11011) );
  CMXI2X1 U20964 ( .A0(n10980), .A1(n11011), .S(n3417), .Z(N5651) );
  CMX2X1 U20965 ( .A0(N7771), .A1(N7770), .S(n4251), .Z(n10987) );
  CMXI2X1 U20966 ( .A0(n10987), .A1(n10981), .S(n4107), .Z(n10994) );
  CMX2X1 U20967 ( .A0(n10982), .A1(n10994), .S(n3772), .Z(n11014) );
  CMXI2X1 U20968 ( .A0(n10983), .A1(n11014), .S(n3417), .Z(N5652) );
  CMX2X1 U20969 ( .A0(N7770), .A1(N7769), .S(n4251), .Z(n10990) );
  CMXI2X1 U20970 ( .A0(n10990), .A1(n10984), .S(n4107), .Z(n10997) );
  CMX2X1 U20971 ( .A0(n10985), .A1(n10997), .S(n3773), .Z(n11017) );
  CMXI2X1 U20972 ( .A0(n10986), .A1(n11017), .S(n3417), .Z(N5653) );
  CMX2X1 U20973 ( .A0(N7769), .A1(N7768), .S(n4251), .Z(n10993) );
  CMXI2X1 U20974 ( .A0(n10993), .A1(n10987), .S(n4107), .Z(n11007) );
  CMX2X1 U20975 ( .A0(n10988), .A1(n11007), .S(n3774), .Z(n11020) );
  CMXI2X1 U20976 ( .A0(n10989), .A1(n11020), .S(n3417), .Z(N5654) );
  CMX2X1 U20977 ( .A0(N7768), .A1(N7767), .S(n4251), .Z(n10996) );
  CMXI2X1 U20978 ( .A0(n10996), .A1(n10990), .S(n4107), .Z(n11010) );
  CMX2X1 U20979 ( .A0(n10991), .A1(n11010), .S(n3775), .Z(n11023) );
  CMXI2X1 U20980 ( .A0(n10992), .A1(n11023), .S(n3420), .Z(N5655) );
  CMX2X1 U20981 ( .A0(N7767), .A1(N7766), .S(n4251), .Z(n11006) );
  CMXI2X1 U20982 ( .A0(n11006), .A1(n10993), .S(n4107), .Z(n11013) );
  CMX2X1 U20983 ( .A0(n10994), .A1(n11013), .S(n3776), .Z(n11026) );
  CMXI2X1 U20984 ( .A0(n10995), .A1(n11026), .S(n3420), .Z(N5656) );
  CMX2X1 U20985 ( .A0(N7766), .A1(N7765), .S(n4251), .Z(n11009) );
  CMXI2X1 U20986 ( .A0(n11009), .A1(n10996), .S(n4107), .Z(n11016) );
  CMX2X1 U20987 ( .A0(n10997), .A1(n11016), .S(n3777), .Z(n11029) );
  CMXI2X1 U20988 ( .A0(n10998), .A1(n11029), .S(n3420), .Z(N5657) );
  CMXI2X1 U20989 ( .A0(n11069), .A1(n10999), .S(n4107), .Z(n11136) );
  CMX2X1 U20990 ( .A0(n11000), .A1(n11136), .S(n3790), .Z(n11269) );
  CMXI2X1 U20991 ( .A0(n11001), .A1(n11269), .S(n3420), .Z(N5207) );
  CMXI2X1 U20992 ( .A0(n4420), .A1(n11003), .S(n3800), .Z(n11005) );
  CMXI2X1 U20993 ( .A0(n11005), .A1(n11004), .S(n3420), .Z(N5162) );
  CMX2X1 U20994 ( .A0(N7765), .A1(N7764), .S(n4251), .Z(n11012) );
  CMXI2X1 U20995 ( .A0(n11012), .A1(n11006), .S(n4107), .Z(n11019) );
  CMX2X1 U20996 ( .A0(n11007), .A1(n11019), .S(n3791), .Z(n11032) );
  CMXI2X1 U20997 ( .A0(n11008), .A1(n11032), .S(n3419), .Z(N5658) );
  CMX2X1 U20998 ( .A0(N7764), .A1(N7763), .S(n4251), .Z(n11015) );
  CMXI2X1 U20999 ( .A0(n11015), .A1(n11009), .S(n4107), .Z(n11022) );
  CMX2X1 U21000 ( .A0(n11010), .A1(n11022), .S(n3797), .Z(n11035) );
  CMXI2X1 U21001 ( .A0(n11011), .A1(n11035), .S(n3419), .Z(N5659) );
  CMX2X1 U21002 ( .A0(N7763), .A1(N7762), .S(n4251), .Z(n11018) );
  CMXI2X1 U21003 ( .A0(n11018), .A1(n11012), .S(n4107), .Z(n11025) );
  CMX2X1 U21004 ( .A0(n11013), .A1(n11025), .S(n3805), .Z(n11041) );
  CMXI2X1 U21005 ( .A0(n11014), .A1(n11041), .S(n3419), .Z(N5660) );
  CMX2X1 U21006 ( .A0(N7762), .A1(N7761), .S(n4251), .Z(n11021) );
  CMXI2X1 U21007 ( .A0(n11021), .A1(n11015), .S(n4107), .Z(n11028) );
  CMX2X1 U21008 ( .A0(n11016), .A1(n11028), .S(n3796), .Z(n11044) );
  CMXI2X1 U21009 ( .A0(n11017), .A1(n11044), .S(n3419), .Z(N5661) );
  CMX2X1 U21010 ( .A0(N7761), .A1(N7760), .S(n4250), .Z(n11024) );
  CMXI2X1 U21011 ( .A0(n11024), .A1(n11018), .S(n4106), .Z(n11031) );
  CMX2X1 U21012 ( .A0(n11019), .A1(n11031), .S(n3797), .Z(n11047) );
  CMXI2X1 U21013 ( .A0(n11020), .A1(n11047), .S(n3419), .Z(N5662) );
  CMX2X1 U21014 ( .A0(N7760), .A1(N7759), .S(n4250), .Z(n11027) );
  CMXI2X1 U21015 ( .A0(n11027), .A1(n11021), .S(n4106), .Z(n11034) );
  CMX2X1 U21016 ( .A0(n11022), .A1(n11034), .S(n3805), .Z(n11050) );
  CMXI2X1 U21017 ( .A0(n11023), .A1(n11050), .S(n3419), .Z(N5663) );
  CMX2X1 U21018 ( .A0(N7759), .A1(N7758), .S(n4250), .Z(n11030) );
  CMXI2X1 U21019 ( .A0(n11030), .A1(n11024), .S(n4106), .Z(n11040) );
  CMX2X1 U21020 ( .A0(n11025), .A1(n11040), .S(n3806), .Z(n11053) );
  CMXI2X1 U21021 ( .A0(n11026), .A1(n11053), .S(n3419), .Z(N5664) );
  CMX2X1 U21022 ( .A0(N7758), .A1(N7757), .S(n4250), .Z(n11033) );
  CMXI2X1 U21023 ( .A0(n11033), .A1(n11027), .S(n4106), .Z(n11043) );
  CMX2X1 U21024 ( .A0(n11028), .A1(n11043), .S(n3807), .Z(n11056) );
  CMXI2X1 U21025 ( .A0(n11029), .A1(n11056), .S(n3419), .Z(N5665) );
  CMX2X1 U21026 ( .A0(N7757), .A1(N7756), .S(n4250), .Z(n11039) );
  CMXI2X1 U21027 ( .A0(n11039), .A1(n11030), .S(n4106), .Z(n11046) );
  CMX2X1 U21028 ( .A0(n11031), .A1(n11046), .S(n3775), .Z(n11059) );
  CMXI2X1 U21029 ( .A0(n11032), .A1(n11059), .S(n3419), .Z(N5666) );
  CMXI2X1 U21030 ( .A0(n11042), .A1(n11033), .S(n4106), .Z(n11049) );
  CMX2X1 U21031 ( .A0(n11034), .A1(n11049), .S(n3792), .Z(n11062) );
  CMXI2X1 U21032 ( .A0(n11035), .A1(n11062), .S(n3419), .Z(N5667) );
  CMX2X1 U21033 ( .A0(N8215), .A1(N8214), .S(n4250), .Z(n11102) );
  CMXI2X1 U21034 ( .A0(n11102), .A1(n11036), .S(n4106), .Z(n11169) );
  CMX2X1 U21035 ( .A0(n11037), .A1(n11169), .S(n3793), .Z(n11302) );
  CMXI2X1 U21036 ( .A0(n11038), .A1(n11302), .S(n3419), .Z(N5208) );
  CMX2X1 U21037 ( .A0(N7755), .A1(N7754), .S(n4250), .Z(n11045) );
  CMXI2X1 U21038 ( .A0(n11045), .A1(n11039), .S(n4106), .Z(n11052) );
  CMX2X1 U21039 ( .A0(n11040), .A1(n11052), .S(n3794), .Z(n11065) );
  CMXI2X1 U21040 ( .A0(n11041), .A1(n11065), .S(n3418), .Z(N5668) );
  CMX2X1 U21041 ( .A0(N7754), .A1(N7753), .S(n4250), .Z(n11048) );
  CMXI2X1 U21042 ( .A0(n11048), .A1(n11042), .S(n4106), .Z(n11055) );
  CMX2X1 U21043 ( .A0(n11043), .A1(n11055), .S(n3795), .Z(n11068) );
  CMXI2X1 U21044 ( .A0(n11044), .A1(n11068), .S(n3418), .Z(N5669) );
  CMX2X1 U21045 ( .A0(N7753), .A1(N7752), .S(n4279), .Z(n11051) );
  CMXI2X1 U21046 ( .A0(n11051), .A1(n11045), .S(n4106), .Z(n11058) );
  CMX2X1 U21047 ( .A0(n11046), .A1(n11058), .S(n3796), .Z(n11074) );
  CMXI2X1 U21048 ( .A0(n11047), .A1(n11074), .S(n3422), .Z(N5670) );
  CMX2X1 U21049 ( .A0(N7752), .A1(N7751), .S(n4261), .Z(n11054) );
  CMXI2X1 U21050 ( .A0(n11054), .A1(n11048), .S(n4106), .Z(n11061) );
  CMX2X1 U21051 ( .A0(n11049), .A1(n11061), .S(n3797), .Z(n11077) );
  CMXI2X1 U21052 ( .A0(n11050), .A1(n11077), .S(n3422), .Z(N5671) );
  CMX2X1 U21053 ( .A0(N7751), .A1(N7750), .S(n3878), .Z(n11057) );
  CMXI2X1 U21054 ( .A0(n11057), .A1(n11051), .S(n4106), .Z(n11064) );
  CMX2X1 U21055 ( .A0(n11052), .A1(n11064), .S(n3805), .Z(n11080) );
  CMXI2X1 U21056 ( .A0(n11053), .A1(n11080), .S(n3421), .Z(N5672) );
  CMX2X1 U21057 ( .A0(N7750), .A1(N7749), .S(n3868), .Z(n11060) );
  CMXI2X1 U21058 ( .A0(n11060), .A1(n11054), .S(n4106), .Z(n11067) );
  CMX2X1 U21059 ( .A0(n11055), .A1(n11067), .S(n3806), .Z(n11083) );
  CMXI2X1 U21060 ( .A0(n11056), .A1(n11083), .S(n3421), .Z(N5673) );
  CMX2X1 U21061 ( .A0(N7749), .A1(N7748), .S(n3869), .Z(n11063) );
  CMXI2X1 U21062 ( .A0(n11063), .A1(n11057), .S(n4106), .Z(n11073) );
  CMX2X1 U21063 ( .A0(n11058), .A1(n11073), .S(n3807), .Z(n11086) );
  CMXI2X1 U21064 ( .A0(n11059), .A1(n11086), .S(n3421), .Z(N5674) );
  CMX2X1 U21065 ( .A0(N7748), .A1(N7747), .S(n3870), .Z(n11066) );
  CMXI2X1 U21066 ( .A0(n11066), .A1(n11060), .S(n4106), .Z(n11076) );
  CMX2X1 U21067 ( .A0(n11061), .A1(n11076), .S(n3808), .Z(n11089) );
  CMXI2X1 U21068 ( .A0(n11062), .A1(n11089), .S(n3421), .Z(N5675) );
  CMX2X1 U21069 ( .A0(N7747), .A1(N7746), .S(n3871), .Z(n11072) );
  CMXI2X1 U21070 ( .A0(n11072), .A1(n11063), .S(n4106), .Z(n11079) );
  CMX2X1 U21071 ( .A0(n11064), .A1(n11079), .S(n3809), .Z(n11092) );
  CMXI2X1 U21072 ( .A0(n11065), .A1(n11092), .S(n3421), .Z(N5676) );
  CMX2X1 U21073 ( .A0(N7746), .A1(N7745), .S(n3867), .Z(n11075) );
  CMXI2X1 U21074 ( .A0(n11075), .A1(n11066), .S(n4105), .Z(n11082) );
  CMX2X1 U21075 ( .A0(n11067), .A1(n11082), .S(n3810), .Z(n11095) );
  CMXI2X1 U21076 ( .A0(n11068), .A1(n11095), .S(n3421), .Z(N5677) );
  CMX2X1 U21077 ( .A0(N8214), .A1(N8213), .S(n3863), .Z(n11135) );
  CMXI2X1 U21078 ( .A0(n11135), .A1(n11069), .S(n4105), .Z(n11202) );
  CMX2X1 U21079 ( .A0(n11070), .A1(n11202), .S(n3811), .Z(n11335) );
  CMXI2X1 U21080 ( .A0(n11071), .A1(n11335), .S(n3421), .Z(N5209) );
  CMX2X1 U21081 ( .A0(N7745), .A1(N7744), .S(n3864), .Z(n11078) );
  CMXI2X1 U21082 ( .A0(n11078), .A1(n11072), .S(n4105), .Z(n11085) );
  CMX2X1 U21083 ( .A0(n11073), .A1(n11085), .S(n3812), .Z(n11098) );
  CMXI2X1 U21084 ( .A0(n11074), .A1(n11098), .S(n3421), .Z(N5678) );
  CMX2X1 U21085 ( .A0(N7744), .A1(N7743), .S(n3865), .Z(n11081) );
  CMXI2X1 U21086 ( .A0(n11081), .A1(n11075), .S(n4105), .Z(n11088) );
  CMX2X1 U21087 ( .A0(n11076), .A1(n11088), .S(n4339), .Z(n11101) );
  CMXI2X1 U21088 ( .A0(n11077), .A1(n11101), .S(n3421), .Z(N5679) );
  CMX2X1 U21089 ( .A0(N7743), .A1(N7742), .S(n3866), .Z(n11084) );
  CMXI2X1 U21090 ( .A0(n11084), .A1(n11078), .S(n4105), .Z(n11091) );
  CMX2X1 U21091 ( .A0(n11079), .A1(n11091), .S(n3771), .Z(n11107) );
  CMXI2X1 U21092 ( .A0(n11080), .A1(n11107), .S(n3421), .Z(N5680) );
  CMX2X1 U21093 ( .A0(N7742), .A1(N7741), .S(n3867), .Z(n11087) );
  CMXI2X1 U21094 ( .A0(n11087), .A1(n11081), .S(n4105), .Z(n11094) );
  CMX2X1 U21095 ( .A0(n11082), .A1(n11094), .S(n3795), .Z(n11110) );
  CMXI2X1 U21096 ( .A0(n11083), .A1(n11110), .S(n3421), .Z(N5681) );
  CMX2X1 U21097 ( .A0(N7741), .A1(N7740), .S(n3868), .Z(n11090) );
  CMXI2X1 U21098 ( .A0(n11090), .A1(n11084), .S(n4105), .Z(n11097) );
  CMX2X1 U21099 ( .A0(n11085), .A1(n11097), .S(n3811), .Z(n11113) );
  CMXI2X1 U21100 ( .A0(n11086), .A1(n11113), .S(n3420), .Z(N5682) );
  CMX2X1 U21101 ( .A0(N7740), .A1(N7739), .S(n3869), .Z(n11093) );
  CMXI2X1 U21102 ( .A0(n11093), .A1(n11087), .S(n4105), .Z(n11100) );
  CMX2X1 U21103 ( .A0(n11088), .A1(n11100), .S(n3797), .Z(n11116) );
  CMXI2X1 U21104 ( .A0(n11089), .A1(n11116), .S(n3420), .Z(N5683) );
  CMX2X1 U21105 ( .A0(N7739), .A1(N7738), .S(n3874), .Z(n11096) );
  CMXI2X1 U21106 ( .A0(n11096), .A1(n11090), .S(n4105), .Z(n11106) );
  CMX2X1 U21107 ( .A0(n11091), .A1(n11106), .S(n3771), .Z(n11119) );
  CMXI2X1 U21108 ( .A0(n11092), .A1(n11119), .S(n3420), .Z(N5684) );
  CMX2X1 U21109 ( .A0(N7738), .A1(N7737), .S(n3875), .Z(n11099) );
  CMXI2X1 U21110 ( .A0(n11099), .A1(n11093), .S(n4105), .Z(n11109) );
  CMX2X1 U21111 ( .A0(n11094), .A1(n11109), .S(n3775), .Z(n11122) );
  CMXI2X1 U21112 ( .A0(n11095), .A1(n11122), .S(n3420), .Z(N5685) );
  CMX2X1 U21113 ( .A0(N7737), .A1(N7736), .S(n3870), .Z(n11105) );
  CMXI2X1 U21114 ( .A0(n11105), .A1(n11096), .S(n4105), .Z(n11112) );
  CMX2X1 U21115 ( .A0(n11097), .A1(n11112), .S(n3811), .Z(n11125) );
  CMXI2X1 U21116 ( .A0(n11098), .A1(n11125), .S(n3420), .Z(N5686) );
  CMX2X1 U21117 ( .A0(N7736), .A1(N7735), .S(n3871), .Z(n11108) );
  CMXI2X1 U21118 ( .A0(n11108), .A1(n11099), .S(n4105), .Z(n11115) );
  CMX2X1 U21119 ( .A0(n11100), .A1(n11115), .S(n3776), .Z(n11128) );
  CMXI2X1 U21120 ( .A0(n11101), .A1(n11128), .S(n3423), .Z(N5687) );
  CMX2X1 U21121 ( .A0(N8213), .A1(N8212), .S(n3872), .Z(n11168) );
  CMXI2X1 U21122 ( .A0(n11168), .A1(n11102), .S(n4105), .Z(n11235) );
  CMX2X1 U21123 ( .A0(n11103), .A1(n11235), .S(n3777), .Z(n11372) );
  CMXI2X1 U21124 ( .A0(n11104), .A1(n11372), .S(n3423), .Z(N5210) );
  CMX2X1 U21125 ( .A0(N7735), .A1(N7734), .S(n3873), .Z(n11111) );
  CMXI2X1 U21126 ( .A0(n11111), .A1(n11105), .S(n4105), .Z(n11118) );
  CMX2X1 U21127 ( .A0(n11106), .A1(n11118), .S(n3790), .Z(n11131) );
  CMXI2X1 U21128 ( .A0(n11107), .A1(n11131), .S(n3423), .Z(N5688) );
  CMX2X1 U21129 ( .A0(N7734), .A1(N7733), .S(n3874), .Z(n11114) );
  CMXI2X1 U21130 ( .A0(n11114), .A1(n11108), .S(n4105), .Z(n11121) );
  CMX2X1 U21131 ( .A0(n11109), .A1(n11121), .S(n3791), .Z(n11134) );
  CMXI2X1 U21132 ( .A0(n11110), .A1(n11134), .S(n3300), .Z(N5689) );
  CMX2X1 U21133 ( .A0(N7733), .A1(N7732), .S(n3875), .Z(n11117) );
  CMXI2X1 U21134 ( .A0(n11117), .A1(n11111), .S(n4105), .Z(n11124) );
  CMX2X1 U21135 ( .A0(n11112), .A1(n11124), .S(n3792), .Z(n11140) );
  CMXI2X1 U21136 ( .A0(n11113), .A1(n11140), .S(n3451), .Z(N5690) );
  CMX2X1 U21137 ( .A0(N7732), .A1(N7731), .S(n3872), .Z(n11120) );
  CMXI2X1 U21138 ( .A0(n11120), .A1(n11114), .S(n4104), .Z(n11127) );
  CMX2X1 U21139 ( .A0(n11115), .A1(n11127), .S(n3811), .Z(n11143) );
  CMXI2X1 U21140 ( .A0(n11116), .A1(n11143), .S(n3429), .Z(N5691) );
  CMX2X1 U21141 ( .A0(N7731), .A1(N7730), .S(n3873), .Z(n11123) );
  CMXI2X1 U21142 ( .A0(n11123), .A1(n11117), .S(n4104), .Z(n11130) );
  CMX2X1 U21143 ( .A0(n11118), .A1(n11130), .S(n3772), .Z(n11146) );
  CMXI2X1 U21144 ( .A0(n11119), .A1(n11146), .S(n3456), .Z(N5692) );
  CMX2X1 U21145 ( .A0(N7730), .A1(N7729), .S(n3874), .Z(n11126) );
  CMXI2X1 U21146 ( .A0(n11126), .A1(n11120), .S(n4104), .Z(n11133) );
  CMX2X1 U21147 ( .A0(n11121), .A1(n11133), .S(n3774), .Z(n11149) );
  CMXI2X1 U21148 ( .A0(n11122), .A1(n11149), .S(n3456), .Z(N5693) );
  CMX2X1 U21149 ( .A0(N7729), .A1(N7728), .S(n3875), .Z(n11129) );
  CMXI2X1 U21150 ( .A0(n11129), .A1(n11123), .S(n4104), .Z(n11139) );
  CMX2X1 U21151 ( .A0(n11124), .A1(n11139), .S(n3775), .Z(n11152) );
  CMXI2X1 U21152 ( .A0(n11125), .A1(n11152), .S(n3456), .Z(N5694) );
  CMX2X1 U21153 ( .A0(N7728), .A1(N7727), .S(n3868), .Z(n11132) );
  CMXI2X1 U21154 ( .A0(n11132), .A1(n11126), .S(n4104), .Z(n11142) );
  CMX2X1 U21155 ( .A0(n11127), .A1(n11142), .S(n3776), .Z(n11155) );
  CMXI2X1 U21156 ( .A0(n11128), .A1(n11155), .S(n3456), .Z(N5695) );
  CMX2X1 U21157 ( .A0(N7727), .A1(N7726), .S(n3872), .Z(n11138) );
  CMXI2X1 U21158 ( .A0(n11138), .A1(n11129), .S(n4104), .Z(n11145) );
  CMX2X1 U21159 ( .A0(n11130), .A1(n11145), .S(n3777), .Z(n11158) );
  CMXI2X1 U21160 ( .A0(n11131), .A1(n11158), .S(n3456), .Z(N5696) );
  CMX2X1 U21161 ( .A0(N7726), .A1(N7725), .S(n3873), .Z(n11141) );
  CMXI2X1 U21162 ( .A0(n11141), .A1(n11132), .S(n4104), .Z(n11148) );
  CMX2X1 U21163 ( .A0(n11133), .A1(n11148), .S(n3790), .Z(n11161) );
  CMXI2X1 U21164 ( .A0(n11134), .A1(n11161), .S(n3456), .Z(N5697) );
  CMX2X1 U21165 ( .A0(N8212), .A1(N8211), .S(n3874), .Z(n11201) );
  CMXI2X1 U21166 ( .A0(n11201), .A1(n11135), .S(n4104), .Z(n11268) );
  CMX2X1 U21167 ( .A0(n11136), .A1(n11268), .S(n3791), .Z(n11405) );
  CMXI2X1 U21168 ( .A0(n11137), .A1(n11405), .S(n3456), .Z(N5211) );
  CMX2X1 U21169 ( .A0(N7725), .A1(N7724), .S(n3875), .Z(n11144) );
  CMXI2X1 U21170 ( .A0(n11144), .A1(n11138), .S(n4104), .Z(n11151) );
  CMX2X1 U21171 ( .A0(n11139), .A1(n11151), .S(n3792), .Z(n11164) );
  CMXI2X1 U21172 ( .A0(n11140), .A1(n11164), .S(n3455), .Z(N5698) );
  CMX2X1 U21173 ( .A0(N7724), .A1(N7723), .S(n3876), .Z(n11147) );
  CMXI2X1 U21174 ( .A0(n11147), .A1(n11141), .S(n4104), .Z(n11154) );
  CMX2X1 U21175 ( .A0(n11142), .A1(n11154), .S(n3793), .Z(n11167) );
  CMXI2X1 U21176 ( .A0(n11143), .A1(n11167), .S(n3455), .Z(N5699) );
  CMX2X1 U21177 ( .A0(N7723), .A1(N7722), .S(n3877), .Z(n11150) );
  CMXI2X1 U21178 ( .A0(n11150), .A1(n11144), .S(n4104), .Z(n11157) );
  CMX2X1 U21179 ( .A0(n11145), .A1(n11157), .S(n3794), .Z(n11173) );
  CMXI2X1 U21180 ( .A0(n11146), .A1(n11173), .S(n3455), .Z(N5700) );
  CMX2X1 U21181 ( .A0(N7722), .A1(N7721), .S(n3878), .Z(n11153) );
  CMXI2X1 U21182 ( .A0(n11153), .A1(n11147), .S(n4104), .Z(n11160) );
  CMX2X1 U21183 ( .A0(n11148), .A1(n11160), .S(n3795), .Z(n11176) );
  CMXI2X1 U21184 ( .A0(n11149), .A1(n11176), .S(n3455), .Z(N5701) );
  CMX2X1 U21185 ( .A0(N7721), .A1(N7720), .S(n3876), .Z(n11156) );
  CMXI2X1 U21186 ( .A0(n11156), .A1(n11150), .S(n4104), .Z(n11163) );
  CMX2X1 U21187 ( .A0(n11151), .A1(n11163), .S(n3796), .Z(n11179) );
  CMXI2X1 U21188 ( .A0(n11152), .A1(n11179), .S(n3455), .Z(N5702) );
  CMX2X1 U21189 ( .A0(N7720), .A1(N7719), .S(n3877), .Z(n11159) );
  CMXI2X1 U21190 ( .A0(n11159), .A1(n11153), .S(n4104), .Z(n11166) );
  CMX2X1 U21191 ( .A0(n11154), .A1(n11166), .S(n3797), .Z(n11182) );
  CMXI2X1 U21192 ( .A0(n11155), .A1(n11182), .S(n3455), .Z(N5703) );
  CMX2X1 U21193 ( .A0(N7719), .A1(N7718), .S(n3879), .Z(n11162) );
  CMXI2X1 U21194 ( .A0(n11162), .A1(n11156), .S(n4104), .Z(n11172) );
  CMX2X1 U21195 ( .A0(n11157), .A1(n11172), .S(n3805), .Z(n11185) );
  CMXI2X1 U21196 ( .A0(n11158), .A1(n11185), .S(n3455), .Z(N5704) );
  CMX2X1 U21197 ( .A0(N7718), .A1(N7717), .S(n3880), .Z(n11165) );
  CMXI2X1 U21198 ( .A0(n11165), .A1(n11159), .S(n4104), .Z(n11175) );
  CMX2X1 U21199 ( .A0(n11160), .A1(n11175), .S(n3806), .Z(n11188) );
  CMXI2X1 U21200 ( .A0(n11161), .A1(n11188), .S(n3455), .Z(N5705) );
  CMX2X1 U21201 ( .A0(N7717), .A1(N7716), .S(n3876), .Z(n11171) );
  CMXI2X1 U21202 ( .A0(n11171), .A1(n11162), .S(n4103), .Z(n11178) );
  CMX2X1 U21203 ( .A0(n11163), .A1(n11178), .S(n3775), .Z(n11191) );
  CMXI2X1 U21204 ( .A0(n11164), .A1(n11191), .S(n3455), .Z(N5706) );
  CMX2X1 U21205 ( .A0(N7716), .A1(N7715), .S(n3877), .Z(n11174) );
  CMXI2X1 U21206 ( .A0(n11174), .A1(n11165), .S(n4103), .Z(n11181) );
  CMX2X1 U21207 ( .A0(n11166), .A1(n11181), .S(n3776), .Z(n11194) );
  CMXI2X1 U21208 ( .A0(n11167), .A1(n11194), .S(n3455), .Z(N5707) );
  CMX2X1 U21209 ( .A0(N8211), .A1(N8210), .S(n3878), .Z(n11234) );
  CMXI2X1 U21210 ( .A0(n11234), .A1(n11168), .S(n4103), .Z(n11301) );
  CMX2X1 U21211 ( .A0(n11169), .A1(n11301), .S(n3794), .Z(n11438) );
  CMXI2X1 U21212 ( .A0(n11170), .A1(n11438), .S(n3454), .Z(N5212) );
  CMX2X1 U21213 ( .A0(N7715), .A1(N7714), .S(n3879), .Z(n11177) );
  CMXI2X1 U21214 ( .A0(n11177), .A1(n11171), .S(n4103), .Z(n11184) );
  CMX2X1 U21215 ( .A0(n11172), .A1(n11184), .S(n3795), .Z(n11197) );
  CMXI2X1 U21216 ( .A0(n11173), .A1(n11197), .S(n3458), .Z(N5708) );
  CMX2X1 U21217 ( .A0(N7714), .A1(N7713), .S(n3876), .Z(n11180) );
  CMXI2X1 U21218 ( .A0(n11180), .A1(n11174), .S(n4103), .Z(n11187) );
  CMX2X1 U21219 ( .A0(n11175), .A1(n11187), .S(n3796), .Z(n11200) );
  CMXI2X1 U21220 ( .A0(n11176), .A1(n11200), .S(n3458), .Z(N5709) );
  CMX2X1 U21221 ( .A0(N7713), .A1(N7712), .S(n3877), .Z(n11183) );
  CMXI2X1 U21222 ( .A0(n11183), .A1(n11177), .S(n4103), .Z(n11190) );
  CMX2X1 U21223 ( .A0(n11178), .A1(n11190), .S(n3797), .Z(n11206) );
  CMXI2X1 U21224 ( .A0(n11179), .A1(n11206), .S(n3458), .Z(N5710) );
  CMX2X1 U21225 ( .A0(N7712), .A1(N7711), .S(n3878), .Z(n11186) );
  CMXI2X1 U21226 ( .A0(n11186), .A1(n11180), .S(n4103), .Z(n11193) );
  CMX2X1 U21227 ( .A0(n11181), .A1(n11193), .S(n3805), .Z(n11209) );
  CMXI2X1 U21228 ( .A0(n11182), .A1(n11209), .S(n3457), .Z(N5711) );
  CMX2X1 U21229 ( .A0(N7711), .A1(N7710), .S(n3879), .Z(n11189) );
  CMXI2X1 U21230 ( .A0(n11189), .A1(n11183), .S(n4103), .Z(n11196) );
  CMX2X1 U21231 ( .A0(n11184), .A1(n11196), .S(n3808), .Z(n11212) );
  CMXI2X1 U21232 ( .A0(n11185), .A1(n11212), .S(n3457), .Z(N5712) );
  CMX2X1 U21233 ( .A0(N7710), .A1(N7709), .S(n3869), .Z(n11192) );
  CMXI2X1 U21234 ( .A0(n11192), .A1(n11186), .S(n4103), .Z(n11199) );
  CMX2X1 U21235 ( .A0(n11187), .A1(n11199), .S(n3807), .Z(n11215) );
  CMXI2X1 U21236 ( .A0(n11188), .A1(n11215), .S(n3457), .Z(N5713) );
  CMX2X1 U21237 ( .A0(N7709), .A1(N7708), .S(n3881), .Z(n11195) );
  CMXI2X1 U21238 ( .A0(n11195), .A1(n11189), .S(n4103), .Z(n11205) );
  CMX2X1 U21239 ( .A0(n11190), .A1(n11205), .S(n3808), .Z(n11218) );
  CMXI2X1 U21240 ( .A0(n11191), .A1(n11218), .S(n3457), .Z(N5714) );
  CMX2X1 U21241 ( .A0(N7708), .A1(N7707), .S(n3862), .Z(n11198) );
  CMXI2X1 U21242 ( .A0(n11198), .A1(n11192), .S(n4103), .Z(n11208) );
  CMX2X1 U21243 ( .A0(n11193), .A1(n11208), .S(n3809), .Z(n11221) );
  CMXI2X1 U21244 ( .A0(n11194), .A1(n11221), .S(n3457), .Z(N5715) );
  CMX2X1 U21245 ( .A0(N7707), .A1(N7706), .S(n3863), .Z(n11204) );
  CMXI2X1 U21246 ( .A0(n11204), .A1(n11195), .S(n4103), .Z(n11211) );
  CMX2X1 U21247 ( .A0(n11196), .A1(n11211), .S(n3810), .Z(n11224) );
  CMXI2X1 U21248 ( .A0(n11197), .A1(n11224), .S(n3457), .Z(N5716) );
  CMX2X1 U21249 ( .A0(N7706), .A1(N7705), .S(n3864), .Z(n11207) );
  CMXI2X1 U21250 ( .A0(n11207), .A1(n11198), .S(n4103), .Z(n11214) );
  CMX2X1 U21251 ( .A0(n11199), .A1(n11214), .S(n3811), .Z(n11227) );
  CMXI2X1 U21252 ( .A0(n11200), .A1(n11227), .S(n3457), .Z(N5717) );
  CMX2X1 U21253 ( .A0(N8210), .A1(N8209), .S(n3865), .Z(n11267) );
  CMXI2X1 U21254 ( .A0(n11267), .A1(n11201), .S(n4103), .Z(n11334) );
  CMX2X1 U21255 ( .A0(n11202), .A1(n11334), .S(n3812), .Z(n11471) );
  CMXI2X1 U21256 ( .A0(n11203), .A1(n11471), .S(n3457), .Z(N5213) );
  CMX2X1 U21257 ( .A0(N7705), .A1(N7704), .S(n3866), .Z(n11210) );
  CMXI2X1 U21258 ( .A0(n11210), .A1(n11204), .S(n4103), .Z(n11217) );
  CMX2X1 U21259 ( .A0(n11205), .A1(n11217), .S(n4322), .Z(n11230) );
  CMXI2X1 U21260 ( .A0(n11206), .A1(n11230), .S(n3457), .Z(N5718) );
  CMX2X1 U21261 ( .A0(N7704), .A1(N7703), .S(n3867), .Z(n11213) );
  CMXI2X1 U21262 ( .A0(n11213), .A1(n11207), .S(n4103), .Z(n11220) );
  CMX2X1 U21263 ( .A0(n11208), .A1(n11220), .S(n3771), .Z(n11233) );
  CMXI2X1 U21264 ( .A0(n11209), .A1(n11233), .S(n3457), .Z(N5719) );
  CMX2X1 U21265 ( .A0(N7703), .A1(N7702), .S(n3878), .Z(n11216) );
  CMXI2X1 U21266 ( .A0(n11216), .A1(n11210), .S(n4102), .Z(n11223) );
  CMX2X1 U21267 ( .A0(n11211), .A1(n11223), .S(n3772), .Z(n11239) );
  CMXI2X1 U21268 ( .A0(n11212), .A1(n11239), .S(n3457), .Z(N5720) );
  CMX2X1 U21269 ( .A0(N7702), .A1(N7701), .S(n3879), .Z(n11219) );
  CMXI2X1 U21270 ( .A0(n11219), .A1(n11213), .S(n4102), .Z(n11226) );
  CMX2X1 U21271 ( .A0(n11214), .A1(n11226), .S(n3773), .Z(n11242) );
  CMXI2X1 U21272 ( .A0(n11215), .A1(n11242), .S(n3456), .Z(N5721) );
  CMX2X1 U21273 ( .A0(N7701), .A1(N7700), .S(n3868), .Z(n11222) );
  CMXI2X1 U21274 ( .A0(n11222), .A1(n11216), .S(n4102), .Z(n11229) );
  CMX2X1 U21275 ( .A0(n11217), .A1(n11229), .S(n3774), .Z(n11245) );
  CMXI2X1 U21276 ( .A0(n11218), .A1(n11245), .S(n3456), .Z(N5722) );
  CMX2X1 U21277 ( .A0(N7700), .A1(N7699), .S(n3869), .Z(n11225) );
  CMXI2X1 U21278 ( .A0(n11225), .A1(n11219), .S(n4102), .Z(n11232) );
  CMX2X1 U21279 ( .A0(n11220), .A1(n11232), .S(n3775), .Z(n11248) );
  CMXI2X1 U21280 ( .A0(n11221), .A1(n11248), .S(n3456), .Z(N5723) );
  CMX2X1 U21281 ( .A0(N7699), .A1(N7698), .S(n3880), .Z(n11228) );
  CMXI2X1 U21282 ( .A0(n11228), .A1(n11222), .S(n4102), .Z(n11238) );
  CMX2X1 U21283 ( .A0(n11223), .A1(n11238), .S(n3776), .Z(n11251) );
  CMXI2X1 U21284 ( .A0(n11224), .A1(n11251), .S(n3456), .Z(N5724) );
  CMX2X1 U21285 ( .A0(N7698), .A1(N7697), .S(n3881), .Z(n11231) );
  CMXI2X1 U21286 ( .A0(n11231), .A1(n11225), .S(n4102), .Z(n11241) );
  CMX2X1 U21287 ( .A0(n11226), .A1(n11241), .S(n3777), .Z(n11254) );
  CMXI2X1 U21288 ( .A0(n11227), .A1(n11254), .S(n3459), .Z(N5725) );
  CMX2X1 U21289 ( .A0(N7697), .A1(N7696), .S(n3862), .Z(n11237) );
  CMXI2X1 U21290 ( .A0(n11237), .A1(n11228), .S(n4102), .Z(n11244) );
  CMX2X1 U21291 ( .A0(n11229), .A1(n11244), .S(n3790), .Z(n11257) );
  CMXI2X1 U21292 ( .A0(n11230), .A1(n11257), .S(n3459), .Z(N5726) );
  CMX2X1 U21293 ( .A0(N7696), .A1(N7695), .S(n3863), .Z(n11240) );
  CMXI2X1 U21294 ( .A0(n11240), .A1(n11231), .S(n4102), .Z(n11247) );
  CMX2X1 U21295 ( .A0(n11232), .A1(n11247), .S(n3791), .Z(n11260) );
  CMXI2X1 U21296 ( .A0(n11233), .A1(n11260), .S(n3459), .Z(N5727) );
  CMX2X1 U21297 ( .A0(N8209), .A1(N8208), .S(n3880), .Z(n11300) );
  CMXI2X1 U21298 ( .A0(n11300), .A1(n11234), .S(n4102), .Z(n11371) );
  CMX2X1 U21299 ( .A0(n11235), .A1(n11371), .S(n3776), .Z(n11504) );
  CMXI2X1 U21300 ( .A0(n11236), .A1(n11504), .S(n3459), .Z(N5214) );
  CMX2X1 U21301 ( .A0(N7695), .A1(N7694), .S(n3881), .Z(n11243) );
  CMXI2X1 U21302 ( .A0(n11243), .A1(n11237), .S(n4102), .Z(n11250) );
  CMX2X1 U21303 ( .A0(n11238), .A1(n11250), .S(n3777), .Z(n11263) );
  CMXI2X1 U21304 ( .A0(n11239), .A1(n11263), .S(n3459), .Z(N5728) );
  CMX2X1 U21305 ( .A0(N7694), .A1(N7693), .S(n3862), .Z(n11246) );
  CMXI2X1 U21306 ( .A0(n11246), .A1(n11240), .S(n4102), .Z(n11253) );
  CMX2X1 U21307 ( .A0(n11241), .A1(n11253), .S(n3806), .Z(n11266) );
  CMXI2X1 U21308 ( .A0(n11242), .A1(n11266), .S(n3459), .Z(N5729) );
  CMX2X1 U21309 ( .A0(N7693), .A1(N7692), .S(n3863), .Z(n11249) );
  CMXI2X1 U21310 ( .A0(n11249), .A1(n11243), .S(n4102), .Z(n11256) );
  CMX2X1 U21311 ( .A0(n11244), .A1(n11256), .S(n3807), .Z(n11272) );
  CMXI2X1 U21312 ( .A0(n11245), .A1(n11272), .S(n3459), .Z(N5730) );
  CMXI2X1 U21313 ( .A0(n11252), .A1(n11246), .S(n4102), .Z(n11259) );
  CMX2X1 U21314 ( .A0(n11247), .A1(n11259), .S(n3808), .Z(n11275) );
  CMXI2X1 U21315 ( .A0(n11248), .A1(n11275), .S(n3459), .Z(N5731) );
  CMX2X1 U21316 ( .A0(N7691), .A1(N7690), .S(n3870), .Z(n11255) );
  CMXI2X1 U21317 ( .A0(n11255), .A1(n11249), .S(n4102), .Z(n11262) );
  CMX2X1 U21318 ( .A0(n11250), .A1(n11262), .S(n3809), .Z(n11278) );
  CMXI2X1 U21319 ( .A0(n11251), .A1(n11278), .S(n3459), .Z(N5732) );
  CMX2X1 U21320 ( .A0(N7690), .A1(N7689), .S(n3871), .Z(n11258) );
  CMXI2X1 U21321 ( .A0(n11258), .A1(n11252), .S(n4102), .Z(n11265) );
  CMX2X1 U21322 ( .A0(n11253), .A1(n11265), .S(n3810), .Z(n11281) );
  CMXI2X1 U21323 ( .A0(n11254), .A1(n11281), .S(n3459), .Z(N5733) );
  CMX2X1 U21324 ( .A0(N7689), .A1(N7688), .S(n3872), .Z(n11261) );
  CMXI2X1 U21325 ( .A0(n11261), .A1(n11255), .S(n4102), .Z(n11271) );
  CMX2X1 U21326 ( .A0(n11256), .A1(n11271), .S(n3809), .Z(n11284) );
  CMXI2X1 U21327 ( .A0(n11257), .A1(n11284), .S(n3458), .Z(N5734) );
  CMX2X1 U21328 ( .A0(N7688), .A1(N7687), .S(n3873), .Z(n11264) );
  CMXI2X1 U21329 ( .A0(n11264), .A1(n11258), .S(n4101), .Z(n11274) );
  CMX2X1 U21330 ( .A0(n11259), .A1(n11274), .S(n3792), .Z(n11287) );
  CMXI2X1 U21331 ( .A0(n11260), .A1(n11287), .S(n3458), .Z(N5735) );
  CMX2X1 U21332 ( .A0(N7687), .A1(N7686), .S(n3874), .Z(n11270) );
  CMXI2X1 U21333 ( .A0(n11270), .A1(n11261), .S(n4101), .Z(n11277) );
  CMX2X1 U21334 ( .A0(n11262), .A1(n11277), .S(n3793), .Z(n11290) );
  CMXI2X1 U21335 ( .A0(n11263), .A1(n11290), .S(n3458), .Z(N5736) );
  CMX2X1 U21336 ( .A0(N7686), .A1(N7685), .S(n3875), .Z(n11273) );
  CMXI2X1 U21337 ( .A0(n11273), .A1(n11264), .S(n4101), .Z(n11280) );
  CMX2X1 U21338 ( .A0(n11265), .A1(n11280), .S(n3794), .Z(n11293) );
  CMXI2X1 U21339 ( .A0(n11266), .A1(n11293), .S(n3458), .Z(N5737) );
  CMX2X1 U21340 ( .A0(N8208), .A1(N8207), .S(n3876), .Z(n11333) );
  CMXI2X1 U21341 ( .A0(n11333), .A1(n11267), .S(n4101), .Z(n11404) );
  CMX2X1 U21342 ( .A0(n11268), .A1(n11404), .S(n3795), .Z(n11537) );
  CMXI2X1 U21343 ( .A0(n11269), .A1(n11537), .S(n3458), .Z(N5215) );
  CMX2X1 U21344 ( .A0(N7685), .A1(N7684), .S(n3880), .Z(n11276) );
  CMXI2X1 U21345 ( .A0(n11276), .A1(n11270), .S(n4101), .Z(n11283) );
  CMX2X1 U21346 ( .A0(n11271), .A1(n11283), .S(n3796), .Z(n11296) );
  CMXI2X1 U21347 ( .A0(n11272), .A1(n11296), .S(n3458), .Z(N5738) );
  CMX2X1 U21348 ( .A0(N7684), .A1(N7683), .S(n3881), .Z(n11279) );
  CMXI2X1 U21349 ( .A0(n11279), .A1(n11273), .S(n4101), .Z(n11286) );
  CMX2X1 U21350 ( .A0(n11274), .A1(n11286), .S(n3797), .Z(n11299) );
  CMXI2X1 U21351 ( .A0(n11275), .A1(n11299), .S(n3458), .Z(N5739) );
  CMX2X1 U21352 ( .A0(N7683), .A1(N7682), .S(n3877), .Z(n11282) );
  CMXI2X1 U21353 ( .A0(n11282), .A1(n11276), .S(n4101), .Z(n11289) );
  CMX2X1 U21354 ( .A0(n11277), .A1(n11289), .S(n3805), .Z(n11305) );
  CMXI2X1 U21355 ( .A0(n11278), .A1(n11305), .S(n3458), .Z(N5740) );
  CMX2X1 U21356 ( .A0(N7682), .A1(N7681), .S(n3878), .Z(n11285) );
  CMXI2X1 U21357 ( .A0(n11285), .A1(n11279), .S(n4101), .Z(n11292) );
  CMX2X1 U21358 ( .A0(n11280), .A1(n11292), .S(n3806), .Z(n11308) );
  CMXI2X1 U21359 ( .A0(n11281), .A1(n11308), .S(n3461), .Z(N5741) );
  CMX2X1 U21360 ( .A0(N7681), .A1(N7680), .S(n3864), .Z(n11288) );
  CMXI2X1 U21361 ( .A0(n11288), .A1(n11282), .S(n4101), .Z(n11295) );
  CMX2X1 U21362 ( .A0(n11283), .A1(n11295), .S(n3807), .Z(n11311) );
  CMXI2X1 U21363 ( .A0(n11284), .A1(n11311), .S(n3461), .Z(N5742) );
  CMX2X1 U21364 ( .A0(N7680), .A1(N7679), .S(n3865), .Z(n11291) );
  CMXI2X1 U21365 ( .A0(n11291), .A1(n11285), .S(n4101), .Z(n11298) );
  CMX2X1 U21366 ( .A0(n11286), .A1(n11298), .S(n3808), .Z(n11314) );
  CMXI2X1 U21367 ( .A0(n11287), .A1(n11314), .S(n3461), .Z(N5743) );
  CMX2X1 U21368 ( .A0(N7679), .A1(N7678), .S(n3866), .Z(n11294) );
  CMXI2X1 U21369 ( .A0(n11294), .A1(n11288), .S(n4101), .Z(n11304) );
  CMX2X1 U21370 ( .A0(n11289), .A1(n11304), .S(n3809), .Z(n11317) );
  CMXI2X1 U21371 ( .A0(n11290), .A1(n11317), .S(n3461), .Z(N5744) );
  CMX2X1 U21372 ( .A0(N7678), .A1(N7677), .S(n3867), .Z(n11297) );
  CMXI2X1 U21373 ( .A0(n11297), .A1(n11291), .S(n4101), .Z(n11307) );
  CMX2X1 U21374 ( .A0(n11292), .A1(n11307), .S(n3810), .Z(n11320) );
  CMXI2X1 U21375 ( .A0(n11293), .A1(n11320), .S(n3461), .Z(N5745) );
  CMX2X1 U21376 ( .A0(N7677), .A1(N7676), .S(n3864), .Z(n11303) );
  CMXI2X1 U21377 ( .A0(n11303), .A1(n11294), .S(n4101), .Z(n11310) );
  CMX2X1 U21378 ( .A0(n11295), .A1(n11310), .S(n3811), .Z(n11323) );
  CMXI2X1 U21379 ( .A0(n11296), .A1(n11323), .S(n3461), .Z(N5746) );
  CMX2X1 U21380 ( .A0(N7676), .A1(N7675), .S(n3865), .Z(n11306) );
  CMXI2X1 U21381 ( .A0(n11306), .A1(n11297), .S(n4101), .Z(n11313) );
  CMX2X1 U21382 ( .A0(n11298), .A1(n11313), .S(n3812), .Z(n11326) );
  CMXI2X1 U21383 ( .A0(n11299), .A1(n11326), .S(n3460), .Z(N5747) );
  CMX2X1 U21384 ( .A0(N8207), .A1(N8206), .S(n3866), .Z(n11370) );
  CMXI2X1 U21385 ( .A0(n11370), .A1(n11300), .S(n4101), .Z(n11437) );
  CMX2X1 U21386 ( .A0(n11301), .A1(n11437), .S(n4320), .Z(n11570) );
  CMXI2X1 U21387 ( .A0(n11302), .A1(n11570), .S(n3460), .Z(N5216) );
  CMX2X1 U21388 ( .A0(N7675), .A1(N7674), .S(n3867), .Z(n11309) );
  CMXI2X1 U21389 ( .A0(n11309), .A1(n11303), .S(n4101), .Z(n11316) );
  CMX2X1 U21390 ( .A0(n11304), .A1(n11316), .S(n3771), .Z(n11329) );
  CMXI2X1 U21391 ( .A0(n11305), .A1(n11329), .S(n3460), .Z(N5748) );
  CMX2X1 U21392 ( .A0(N7674), .A1(N7673), .S(n3871), .Z(n11312) );
  CMXI2X1 U21393 ( .A0(n11312), .A1(n11306), .S(n4100), .Z(n11319) );
  CMX2X1 U21394 ( .A0(n11307), .A1(n11319), .S(n3777), .Z(n11332) );
  CMXI2X1 U21395 ( .A0(n11308), .A1(n11332), .S(n3460), .Z(N5749) );
  CMX2X1 U21396 ( .A0(N7673), .A1(N7672), .S(n3879), .Z(n11315) );
  CMXI2X1 U21397 ( .A0(n11315), .A1(n11309), .S(n4100), .Z(n11322) );
  CMX2X1 U21398 ( .A0(n11310), .A1(n11322), .S(n3790), .Z(n11342) );
  CMXI2X1 U21399 ( .A0(n11311), .A1(n11342), .S(n3460), .Z(N5750) );
  CMX2X1 U21400 ( .A0(N7672), .A1(N7671), .S(n3880), .Z(n11318) );
  CMXI2X1 U21401 ( .A0(n11318), .A1(n11312), .S(n4100), .Z(n11325) );
  CMX2X1 U21402 ( .A0(n11313), .A1(n11325), .S(n3811), .Z(n11345) );
  CMXI2X1 U21403 ( .A0(n11314), .A1(n11345), .S(n3460), .Z(N5751) );
  CMX2X1 U21404 ( .A0(N7671), .A1(N7670), .S(n3881), .Z(n11321) );
  CMXI2X1 U21405 ( .A0(n11321), .A1(n11315), .S(n4100), .Z(n11328) );
  CMX2X1 U21406 ( .A0(n11316), .A1(n11328), .S(n3812), .Z(n11348) );
  CMXI2X1 U21407 ( .A0(n11317), .A1(n11348), .S(n3460), .Z(N5752) );
  CMX2X1 U21408 ( .A0(N7670), .A1(N7669), .S(n3862), .Z(n11324) );
  CMXI2X1 U21409 ( .A0(n11324), .A1(n11318), .S(n4100), .Z(n11331) );
  CMX2X1 U21410 ( .A0(n11319), .A1(n11331), .S(n4314), .Z(n11351) );
  CMXI2X1 U21411 ( .A0(n11320), .A1(n11351), .S(n3460), .Z(N5753) );
  CMX2X1 U21412 ( .A0(N7669), .A1(N7668), .S(n3863), .Z(n11327) );
  CMXI2X1 U21413 ( .A0(n11327), .A1(n11321), .S(n4100), .Z(n11341) );
  CMX2X1 U21414 ( .A0(n11322), .A1(n11341), .S(n3771), .Z(n11354) );
  CMXI2X1 U21415 ( .A0(n11323), .A1(n11354), .S(n3460), .Z(N5754) );
  CMX2X1 U21416 ( .A0(N7668), .A1(N7667), .S(n3864), .Z(n11330) );
  CMXI2X1 U21417 ( .A0(n11330), .A1(n11324), .S(n4100), .Z(n11344) );
  CMX2X1 U21418 ( .A0(n11325), .A1(n11344), .S(n3772), .Z(n11357) );
  CMXI2X1 U21419 ( .A0(n11326), .A1(n11357), .S(n3460), .Z(N5755) );
  CMX2X1 U21420 ( .A0(N7667), .A1(N7666), .S(n3865), .Z(n11340) );
  CMXI2X1 U21421 ( .A0(n11340), .A1(n11327), .S(n4100), .Z(n11347) );
  CMX2X1 U21422 ( .A0(n11328), .A1(n11347), .S(n3810), .Z(n11360) );
  CMXI2X1 U21423 ( .A0(n11329), .A1(n11360), .S(n3460), .Z(N5756) );
  CMX2X1 U21424 ( .A0(N7666), .A1(N7665), .S(n3862), .Z(n11343) );
  CMXI2X1 U21425 ( .A0(n11343), .A1(n11330), .S(n4100), .Z(n11350) );
  CMX2X1 U21426 ( .A0(n11331), .A1(n11350), .S(n3772), .Z(n11363) );
  CMXI2X1 U21427 ( .A0(n11332), .A1(n11363), .S(n3459), .Z(N5757) );
  CMX2X1 U21428 ( .A0(N8206), .A1(N8205), .S(n3863), .Z(n11403) );
  CMXI2X1 U21429 ( .A0(n11403), .A1(n11333), .S(n4100), .Z(n11470) );
  CMX2X1 U21430 ( .A0(n11334), .A1(n11470), .S(n3773), .Z(n11603) );
  CMXI2X1 U21431 ( .A0(n11335), .A1(n11603), .S(n3463), .Z(N5217) );
  CMXI2X1 U21432 ( .A0(n4423), .A1(n11337), .S(n3785), .Z(n11339) );
  CMXI2X1 U21433 ( .A0(n11339), .A1(n11338), .S(n3463), .Z(N5163) );
  CMX2X1 U21434 ( .A0(N7665), .A1(N7664), .S(n3866), .Z(n11346) );
  CMXI2X1 U21435 ( .A0(n11346), .A1(n11340), .S(n4100), .Z(n11353) );
  CMX2X1 U21436 ( .A0(n11341), .A1(n11353), .S(n3774), .Z(n11366) );
  CMXI2X1 U21437 ( .A0(n11342), .A1(n11366), .S(n3462), .Z(N5758) );
  CMX2X1 U21438 ( .A0(N7664), .A1(N7663), .S(n3868), .Z(n11349) );
  CMXI2X1 U21439 ( .A0(n11349), .A1(n11343), .S(n4100), .Z(n11356) );
  CMX2X1 U21440 ( .A0(n11344), .A1(n11356), .S(n3775), .Z(n11369) );
  CMXI2X1 U21441 ( .A0(n11345), .A1(n11369), .S(n3462), .Z(N5759) );
  CMX2X1 U21442 ( .A0(N7663), .A1(N7662), .S(n3869), .Z(n11352) );
  CMXI2X1 U21443 ( .A0(n11352), .A1(n11346), .S(n4100), .Z(n11359) );
  CMX2X1 U21444 ( .A0(n11347), .A1(n11359), .S(n3776), .Z(n11375) );
  CMXI2X1 U21445 ( .A0(n11348), .A1(n11375), .S(n3462), .Z(N5760) );
  CMX2X1 U21446 ( .A0(N7662), .A1(N7661), .S(n3870), .Z(n11355) );
  CMXI2X1 U21447 ( .A0(n11355), .A1(n11349), .S(n4100), .Z(n11362) );
  CMX2X1 U21448 ( .A0(n11350), .A1(n11362), .S(n3777), .Z(n11378) );
  CMXI2X1 U21449 ( .A0(n11351), .A1(n11378), .S(n3462), .Z(N5761) );
  CMX2X1 U21450 ( .A0(N7661), .A1(N7660), .S(n3871), .Z(n11358) );
  CMXI2X1 U21451 ( .A0(n11358), .A1(n11352), .S(n4100), .Z(n11365) );
  CMX2X1 U21452 ( .A0(n11353), .A1(n11365), .S(n3790), .Z(n11381) );
  CMXI2X1 U21453 ( .A0(n11354), .A1(n11381), .S(n3462), .Z(N5762) );
  CMX2X1 U21454 ( .A0(N7660), .A1(N7659), .S(n3868), .Z(n11361) );
  CMXI2X1 U21455 ( .A0(n11361), .A1(n11355), .S(n4100), .Z(n11368) );
  CMX2X1 U21456 ( .A0(n11356), .A1(n11368), .S(n3791), .Z(n11384) );
  CMXI2X1 U21457 ( .A0(n11357), .A1(n11384), .S(n3462), .Z(N5763) );
  CMX2X1 U21458 ( .A0(N7659), .A1(N7658), .S(n3869), .Z(n11364) );
  CMXI2X1 U21459 ( .A0(n11364), .A1(n11358), .S(n4099), .Z(n11374) );
  CMX2X1 U21460 ( .A0(n11359), .A1(n11374), .S(n3792), .Z(n11387) );
  CMXI2X1 U21461 ( .A0(n11360), .A1(n11387), .S(n3462), .Z(N5764) );
  CMX2X1 U21462 ( .A0(N7658), .A1(N7657), .S(n3866), .Z(n11367) );
  CMXI2X1 U21463 ( .A0(n11367), .A1(n11361), .S(n4099), .Z(n11377) );
  CMX2X1 U21464 ( .A0(n11362), .A1(n11377), .S(n3793), .Z(n11390) );
  CMXI2X1 U21465 ( .A0(n11363), .A1(n11390), .S(n3462), .Z(N5765) );
  CMX2X1 U21466 ( .A0(N7657), .A1(N7656), .S(n3867), .Z(n11373) );
  CMXI2X1 U21467 ( .A0(n11373), .A1(n11364), .S(n4099), .Z(n11380) );
  CMX2X1 U21468 ( .A0(n11365), .A1(n11380), .S(n3794), .Z(n11393) );
  CMXI2X1 U21469 ( .A0(n11366), .A1(n11393), .S(n3462), .Z(N5766) );
  CMX2X1 U21470 ( .A0(N7656), .A1(N7655), .S(n3868), .Z(n11376) );
  CMXI2X1 U21471 ( .A0(n11376), .A1(n11367), .S(n4099), .Z(n11383) );
  CMX2X1 U21472 ( .A0(n11368), .A1(n11383), .S(n3795), .Z(n11396) );
  CMXI2X1 U21473 ( .A0(n11369), .A1(n11396), .S(n3462), .Z(N5767) );
  CMX2X1 U21474 ( .A0(N8205), .A1(N8204), .S(n3869), .Z(n11436) );
  CMXI2X1 U21475 ( .A0(n11436), .A1(n11370), .S(n4099), .Z(n11503) );
  CMX2X1 U21476 ( .A0(n11371), .A1(n11503), .S(n3796), .Z(n11636) );
  CMXI2X1 U21477 ( .A0(n11372), .A1(n11636), .S(n3462), .Z(N5218) );
  CMX2X1 U21478 ( .A0(N7655), .A1(N7654), .S(n3870), .Z(n11379) );
  CMXI2X1 U21479 ( .A0(n11379), .A1(n11373), .S(n4099), .Z(n11386) );
  CMX2X1 U21480 ( .A0(n11374), .A1(n11386), .S(n3797), .Z(n11399) );
  CMXI2X1 U21481 ( .A0(n11375), .A1(n11399), .S(n3461), .Z(N5768) );
  CMX2X1 U21482 ( .A0(N7654), .A1(N7653), .S(n3871), .Z(n11382) );
  CMXI2X1 U21483 ( .A0(n11382), .A1(n11376), .S(n4099), .Z(n11389) );
  CMX2X1 U21484 ( .A0(n11377), .A1(n11389), .S(n3805), .Z(n11402) );
  CMXI2X1 U21485 ( .A0(n11378), .A1(n11402), .S(n3461), .Z(N5769) );
  CMX2X1 U21486 ( .A0(N7653), .A1(N7652), .S(n3872), .Z(n11385) );
  CMXI2X1 U21487 ( .A0(n11385), .A1(n11379), .S(n4099), .Z(n11392) );
  CMX2X1 U21488 ( .A0(n11380), .A1(n11392), .S(n3790), .Z(n11408) );
  CMXI2X1 U21489 ( .A0(n11381), .A1(n11408), .S(n3461), .Z(N5770) );
  CMX2X1 U21490 ( .A0(N7652), .A1(N7651), .S(n3873), .Z(n11388) );
  CMXI2X1 U21491 ( .A0(n11388), .A1(n11382), .S(n4099), .Z(n11395) );
  CMX2X1 U21492 ( .A0(n11383), .A1(n11395), .S(n3791), .Z(n11411) );
  CMXI2X1 U21493 ( .A0(n11384), .A1(n11411), .S(n3461), .Z(N5771) );
  CMX2X1 U21494 ( .A0(N7651), .A1(N7650), .S(n3880), .Z(n11391) );
  CMXI2X1 U21495 ( .A0(n11391), .A1(n11385), .S(n4099), .Z(n11398) );
  CMX2X1 U21496 ( .A0(n11386), .A1(n11398), .S(n3776), .Z(n11414) );
  CMXI2X1 U21497 ( .A0(n11387), .A1(n11414), .S(n3461), .Z(N5772) );
  CMX2X1 U21498 ( .A0(N7650), .A1(N7649), .S(n3868), .Z(n11394) );
  CMXI2X1 U21499 ( .A0(n11394), .A1(n11388), .S(n4099), .Z(n11401) );
  CMX2X1 U21500 ( .A0(n11389), .A1(n11401), .S(n3777), .Z(n11417) );
  CMXI2X1 U21501 ( .A0(n11390), .A1(n11417), .S(n3430), .Z(N5773) );
  CMX2X1 U21502 ( .A0(N7649), .A1(N7648), .S(n3869), .Z(n11397) );
  CMXI2X1 U21503 ( .A0(n11397), .A1(n11391), .S(n4099), .Z(n11407) );
  CMX2X1 U21504 ( .A0(n11392), .A1(n11407), .S(n3790), .Z(n11420) );
  CMXI2X1 U21505 ( .A0(n11393), .A1(n11420), .S(n3430), .Z(N5774) );
  CMX2X1 U21506 ( .A0(N7648), .A1(N7647), .S(n3870), .Z(n11400) );
  CMXI2X1 U21507 ( .A0(n11400), .A1(n11394), .S(n4099), .Z(n11410) );
  CMX2X1 U21508 ( .A0(n11395), .A1(n11410), .S(n3791), .Z(n11423) );
  CMXI2X1 U21509 ( .A0(n11396), .A1(n11423), .S(n3430), .Z(N5775) );
  CMX2X1 U21510 ( .A0(N7647), .A1(N7646), .S(n3871), .Z(n11406) );
  CMXI2X1 U21511 ( .A0(n11406), .A1(n11397), .S(n4099), .Z(n11413) );
  CMX2X1 U21512 ( .A0(n11398), .A1(n11413), .S(n3792), .Z(n11426) );
  CMXI2X1 U21513 ( .A0(n11399), .A1(n11426), .S(n3429), .Z(N5776) );
  CMX2X1 U21514 ( .A0(N7646), .A1(N7645), .S(n3872), .Z(n11409) );
  CMXI2X1 U21515 ( .A0(n11409), .A1(n11400), .S(n4099), .Z(n11416) );
  CMX2X1 U21516 ( .A0(n11401), .A1(n11416), .S(n3793), .Z(n11429) );
  CMXI2X1 U21517 ( .A0(n11402), .A1(n11429), .S(n3429), .Z(N5777) );
  CMX2X1 U21518 ( .A0(N8204), .A1(N8203), .S(n3873), .Z(n11469) );
  CMXI2X1 U21519 ( .A0(n11469), .A1(n11403), .S(n4099), .Z(n11536) );
  CMX2X1 U21520 ( .A0(n11404), .A1(n11536), .S(n3794), .Z(n11669) );
  CMXI2X1 U21521 ( .A0(n11405), .A1(n11669), .S(n3429), .Z(N5219) );
  CMX2X1 U21522 ( .A0(N7645), .A1(N7644), .S(n3874), .Z(n11412) );
  CMXI2X1 U21523 ( .A0(n11412), .A1(n11406), .S(n4098), .Z(n11419) );
  CMX2X1 U21524 ( .A0(n11407), .A1(n11419), .S(n3795), .Z(n11432) );
  CMXI2X1 U21525 ( .A0(n11408), .A1(n11432), .S(n3429), .Z(N5778) );
  CMX2X1 U21526 ( .A0(N7644), .A1(N7643), .S(n3864), .Z(n11415) );
  CMXI2X1 U21527 ( .A0(n11415), .A1(n11409), .S(n4098), .Z(n11422) );
  CMX2X1 U21528 ( .A0(n11410), .A1(n11422), .S(n3796), .Z(n11435) );
  CMXI2X1 U21529 ( .A0(n11411), .A1(n11435), .S(n3429), .Z(N5779) );
  CMX2X1 U21530 ( .A0(N7643), .A1(N7642), .S(n3865), .Z(n11418) );
  CMXI2X1 U21531 ( .A0(n11418), .A1(n11412), .S(n4098), .Z(n11425) );
  CMX2X1 U21532 ( .A0(n11413), .A1(n11425), .S(n3797), .Z(n11441) );
  CMXI2X1 U21533 ( .A0(n11414), .A1(n11441), .S(n3429), .Z(N5780) );
  CMX2X1 U21534 ( .A0(N7642), .A1(N7641), .S(n3875), .Z(n11421) );
  CMXI2X1 U21535 ( .A0(n11421), .A1(n11415), .S(n4098), .Z(n11428) );
  CMX2X1 U21536 ( .A0(n11416), .A1(n11428), .S(n3805), .Z(n11444) );
  CMXI2X1 U21537 ( .A0(n11417), .A1(n11444), .S(n3429), .Z(N5781) );
  CMX2X1 U21538 ( .A0(N7641), .A1(N7640), .S(n3876), .Z(n11424) );
  CMXI2X1 U21539 ( .A0(n11424), .A1(n11418), .S(n4098), .Z(n11431) );
  CMX2X1 U21540 ( .A0(n11419), .A1(n11431), .S(n3773), .Z(n11447) );
  CMXI2X1 U21541 ( .A0(n11420), .A1(n11447), .S(n3437), .Z(N5782) );
  CMX2X1 U21542 ( .A0(N7640), .A1(N7639), .S(n3870), .Z(n11427) );
  CMXI2X1 U21543 ( .A0(n11427), .A1(n11421), .S(n4098), .Z(n11434) );
  CMX2X1 U21544 ( .A0(n11422), .A1(n11434), .S(n3774), .Z(n11450) );
  CMXI2X1 U21545 ( .A0(n11423), .A1(n11450), .S(n3463), .Z(N5783) );
  CMX2X1 U21546 ( .A0(N7639), .A1(N7638), .S(n3871), .Z(n11430) );
  CMXI2X1 U21547 ( .A0(n11430), .A1(n11424), .S(n4098), .Z(n11440) );
  CMX2X1 U21548 ( .A0(n11425), .A1(n11440), .S(n3775), .Z(n11453) );
  CMXI2X1 U21549 ( .A0(n11426), .A1(n11453), .S(n3463), .Z(N5784) );
  CMX2X1 U21550 ( .A0(N7638), .A1(N7637), .S(n3870), .Z(n11433) );
  CMXI2X1 U21551 ( .A0(n11433), .A1(n11427), .S(n4098), .Z(n11443) );
  CMX2X1 U21552 ( .A0(n11428), .A1(n11443), .S(n3776), .Z(n11456) );
  CMXI2X1 U21553 ( .A0(n11429), .A1(n11456), .S(n3463), .Z(N5785) );
  CMX2X1 U21554 ( .A0(N7637), .A1(N7636), .S(n3871), .Z(n11439) );
  CMXI2X1 U21555 ( .A0(n11439), .A1(n11430), .S(n4098), .Z(n11446) );
  CMX2X1 U21556 ( .A0(n11431), .A1(n11446), .S(n3777), .Z(n11459) );
  CMXI2X1 U21557 ( .A0(n11432), .A1(n11459), .S(n3463), .Z(N5786) );
  CMX2X1 U21558 ( .A0(N7636), .A1(N7635), .S(n3872), .Z(n11442) );
  CMXI2X1 U21559 ( .A0(n11442), .A1(n11433), .S(n4098), .Z(n11449) );
  CMX2X1 U21560 ( .A0(n11434), .A1(n11449), .S(n3811), .Z(n11462) );
  CMXI2X1 U21561 ( .A0(n11435), .A1(n11462), .S(n3463), .Z(N5787) );
  CMX2X1 U21562 ( .A0(N8203), .A1(N8202), .S(n3868), .Z(n11502) );
  CMXI2X1 U21563 ( .A0(n11502), .A1(n11436), .S(n4098), .Z(n11569) );
  CMX2X1 U21564 ( .A0(n11437), .A1(n11569), .S(n3807), .Z(n11706) );
  CMXI2X1 U21565 ( .A0(n11438), .A1(n11706), .S(n3463), .Z(N5220) );
  CMX2X1 U21566 ( .A0(N7635), .A1(N7634), .S(n3869), .Z(n11445) );
  CMXI2X1 U21567 ( .A0(n11445), .A1(n11439), .S(n4098), .Z(n11452) );
  CMX2X1 U21568 ( .A0(n11440), .A1(n11452), .S(n3808), .Z(n11465) );
  CMXI2X1 U21569 ( .A0(n11441), .A1(n11465), .S(n3431), .Z(N5788) );
  CMX2X1 U21570 ( .A0(N7634), .A1(N7633), .S(n3870), .Z(n11448) );
  CMXI2X1 U21571 ( .A0(n11448), .A1(n11442), .S(n4098), .Z(n11455) );
  CMX2X1 U21572 ( .A0(n11443), .A1(n11455), .S(n3809), .Z(n11468) );
  CMXI2X1 U21573 ( .A0(n11444), .A1(n11468), .S(n3431), .Z(N5789) );
  CMX2X1 U21574 ( .A0(N7633), .A1(N7632), .S(n3871), .Z(n11451) );
  CMXI2X1 U21575 ( .A0(n11451), .A1(n11445), .S(n4098), .Z(n11458) );
  CMX2X1 U21576 ( .A0(n11446), .A1(n11458), .S(n3810), .Z(n11474) );
  CMXI2X1 U21577 ( .A0(n11447), .A1(n11474), .S(n3431), .Z(N5790) );
  CMX2X1 U21578 ( .A0(N7632), .A1(N7631), .S(n3872), .Z(n11454) );
  CMXI2X1 U21579 ( .A0(n11454), .A1(n11448), .S(n4098), .Z(n11461) );
  CMX2X1 U21580 ( .A0(n11449), .A1(n11461), .S(n3811), .Z(n11477) );
  CMXI2X1 U21581 ( .A0(n11450), .A1(n11477), .S(n3431), .Z(N5791) );
  CMX2X1 U21582 ( .A0(N7631), .A1(N7630), .S(n3873), .Z(n11457) );
  CMXI2X1 U21583 ( .A0(n11457), .A1(n11451), .S(n4098), .Z(n11464) );
  CMX2X1 U21584 ( .A0(n11452), .A1(n11464), .S(n3812), .Z(n11480) );
  CMXI2X1 U21585 ( .A0(n11453), .A1(n11480), .S(n3431), .Z(N5792) );
  CMX2X1 U21586 ( .A0(N7630), .A1(N7629), .S(n3874), .Z(n11460) );
  CMXI2X1 U21587 ( .A0(n11460), .A1(n11454), .S(n4097), .Z(n11467) );
  CMX2X1 U21588 ( .A0(n11455), .A1(n11467), .S(n4318), .Z(n11483) );
  CMXI2X1 U21589 ( .A0(n11456), .A1(n11483), .S(n3431), .Z(N5793) );
  CMX2X1 U21590 ( .A0(N7629), .A1(N7628), .S(n3864), .Z(n11463) );
  CMXI2X1 U21591 ( .A0(n11463), .A1(n11457), .S(n4097), .Z(n11473) );
  CMX2X1 U21592 ( .A0(n11458), .A1(n11473), .S(n3771), .Z(n11486) );
  CMXI2X1 U21593 ( .A0(n11459), .A1(n11486), .S(n3431), .Z(N5794) );
  CMXI2X1 U21594 ( .A0(n11466), .A1(n11460), .S(n4097), .Z(n11476) );
  CMX2X1 U21595 ( .A0(n11461), .A1(n11476), .S(n3772), .Z(n11489) );
  CMXI2X1 U21596 ( .A0(n11462), .A1(n11489), .S(n3431), .Z(N5795) );
  CMX2X1 U21597 ( .A0(N7627), .A1(N7626), .S(n3875), .Z(n11472) );
  CMXI2X1 U21598 ( .A0(n11472), .A1(n11463), .S(n4097), .Z(n11479) );
  CMX2X1 U21599 ( .A0(n11464), .A1(n11479), .S(n3773), .Z(n11492) );
  CMXI2X1 U21600 ( .A0(n11465), .A1(n11492), .S(n3431), .Z(N5796) );
  CMX2X1 U21601 ( .A0(N7626), .A1(N7625), .S(n3876), .Z(n11475) );
  CMXI2X1 U21602 ( .A0(n11475), .A1(n11466), .S(n4097), .Z(n11482) );
  CMX2X1 U21603 ( .A0(n11467), .A1(n11482), .S(n3774), .Z(n11495) );
  CMXI2X1 U21604 ( .A0(n11468), .A1(n11495), .S(n3431), .Z(N5797) );
  CMX2X1 U21605 ( .A0(N8202), .A1(N8201), .S(n3872), .Z(n11535) );
  CMXI2X1 U21606 ( .A0(n11535), .A1(n11469), .S(n4097), .Z(n11602) );
  CMX2X1 U21607 ( .A0(n11470), .A1(n11602), .S(n3775), .Z(n11739) );
  CMXI2X1 U21608 ( .A0(n11471), .A1(n11739), .S(n3430), .Z(N5221) );
  CMX2X1 U21609 ( .A0(N7625), .A1(N7624), .S(n3873), .Z(n11478) );
  CMXI2X1 U21610 ( .A0(n11478), .A1(n11472), .S(n4097), .Z(n11485) );
  CMX2X1 U21611 ( .A0(n11473), .A1(n11485), .S(n3776), .Z(n11498) );
  CMXI2X1 U21612 ( .A0(n11474), .A1(n11498), .S(n3430), .Z(N5798) );
  CMX2X1 U21613 ( .A0(N7624), .A1(N7623), .S(n3874), .Z(n11481) );
  CMXI2X1 U21614 ( .A0(n11481), .A1(n11475), .S(n4097), .Z(n11488) );
  CMX2X1 U21615 ( .A0(n11476), .A1(n11488), .S(n3777), .Z(n11501) );
  CMXI2X1 U21616 ( .A0(n11477), .A1(n11501), .S(n3430), .Z(N5799) );
  CMX2X1 U21617 ( .A0(N7623), .A1(N7622), .S(n3875), .Z(n11484) );
  CMXI2X1 U21618 ( .A0(n11484), .A1(n11478), .S(n4097), .Z(n11491) );
  CMX2X1 U21619 ( .A0(n11479), .A1(n11491), .S(n3790), .Z(n11507) );
  CMXI2X1 U21620 ( .A0(n11480), .A1(n11507), .S(n3430), .Z(N5800) );
  CMX2X1 U21621 ( .A0(N7622), .A1(N7621), .S(n3872), .Z(n11487) );
  CMXI2X1 U21622 ( .A0(n11487), .A1(n11481), .S(n4097), .Z(n11494) );
  CMX2X1 U21623 ( .A0(n11482), .A1(n11494), .S(n3791), .Z(n11510) );
  CMX2X1 U21624 ( .A0(N7621), .A1(N7620), .S(n3873), .Z(n11490) );
  CMXI2X1 U21625 ( .A0(n11490), .A1(n11484), .S(n4097), .Z(n11497) );
  CMX2X1 U21626 ( .A0(n11485), .A1(n11497), .S(n3791), .Z(n11513) );
  CMX2X1 U21627 ( .A0(N7620), .A1(N7619), .S(n3874), .Z(n11493) );
  CMXI2X1 U21628 ( .A0(n11493), .A1(n11487), .S(n4097), .Z(n11500) );
  CMX2X1 U21629 ( .A0(n11488), .A1(n11500), .S(n3792), .Z(n11516) );
  CMX2X1 U21630 ( .A0(N7619), .A1(N7618), .S(n3875), .Z(n11496) );
  CMXI2X1 U21631 ( .A0(n11496), .A1(n11490), .S(n4097), .Z(n11506) );
  CMX2X1 U21632 ( .A0(n11491), .A1(n11506), .S(n3790), .Z(n11519) );
  CMXI2X1 U21633 ( .A0(n11492), .A1(n11519), .S(n3430), .Z(N5804) );
  CMX2X1 U21634 ( .A0(N7618), .A1(N7617), .S(n3873), .Z(n11499) );
  CMXI2X1 U21635 ( .A0(n11499), .A1(n11493), .S(n4097), .Z(n11509) );
  CMX2X1 U21636 ( .A0(n11494), .A1(n11509), .S(n3791), .Z(n11522) );
  CMXI2X1 U21637 ( .A0(n11495), .A1(n11522), .S(n3433), .Z(N5805) );
  CMX2X1 U21638 ( .A0(N7617), .A1(N7616), .S(n3877), .Z(n11505) );
  CMXI2X1 U21639 ( .A0(n11505), .A1(n11496), .S(n4097), .Z(n11512) );
  CMX2X1 U21640 ( .A0(n11497), .A1(n11512), .S(n3792), .Z(n11525) );
  CMXI2X1 U21641 ( .A0(n11498), .A1(n11525), .S(n3433), .Z(N5806) );
  CMX2X1 U21642 ( .A0(N7616), .A1(N7615), .S(n3878), .Z(n11508) );
  CMXI2X1 U21643 ( .A0(n11508), .A1(n11499), .S(n4097), .Z(n11515) );
  CMX2X1 U21644 ( .A0(n11500), .A1(n11515), .S(n3793), .Z(n11528) );
  CMXI2X1 U21645 ( .A0(n11501), .A1(n11528), .S(n3433), .Z(N5807) );
  CMX2X1 U21646 ( .A0(N8201), .A1(N8200), .S(n3879), .Z(n11568) );
  CMXI2X1 U21647 ( .A0(n11568), .A1(n11502), .S(n4096), .Z(n11635) );
  CMX2X1 U21648 ( .A0(n11503), .A1(n11635), .S(n3794), .Z(n11772) );
  CMXI2X1 U21649 ( .A0(n11504), .A1(n11772), .S(n3433), .Z(N5222) );
  CMX2X1 U21650 ( .A0(N7615), .A1(N7614), .S(n3880), .Z(n11511) );
  CMXI2X1 U21651 ( .A0(n11511), .A1(n11505), .S(n4096), .Z(n11518) );
  CMX2X1 U21652 ( .A0(n11506), .A1(n11518), .S(n3812), .Z(n11531) );
  CMXI2X1 U21653 ( .A0(n11507), .A1(n11531), .S(n3433), .Z(N5808) );
  CMX2X1 U21654 ( .A0(N7614), .A1(N7613), .S(n3881), .Z(n11514) );
  CMXI2X1 U21655 ( .A0(n11514), .A1(n11508), .S(n4096), .Z(n11521) );
  CMX2X1 U21656 ( .A0(n11509), .A1(n11521), .S(n3792), .Z(n11534) );
  CMXI2X1 U21657 ( .A0(n11510), .A1(n11534), .S(n3433), .Z(N5809) );
  CMX2X1 U21658 ( .A0(N7613), .A1(N7612), .S(n3862), .Z(n11517) );
  CMXI2X1 U21659 ( .A0(n11517), .A1(n11511), .S(n4096), .Z(n11524) );
  CMX2X1 U21660 ( .A0(n11512), .A1(n11524), .S(n3793), .Z(n11540) );
  CMXI2X1 U21661 ( .A0(n11513), .A1(n11540), .S(n3432), .Z(N5810) );
  CMX2X1 U21662 ( .A0(N7612), .A1(N7611), .S(n3863), .Z(n11520) );
  CMXI2X1 U21663 ( .A0(n11520), .A1(n11514), .S(n4096), .Z(n11527) );
  CMX2X1 U21664 ( .A0(n11515), .A1(n11527), .S(n3794), .Z(n11543) );
  CMXI2X1 U21665 ( .A0(n11516), .A1(n11543), .S(n3432), .Z(N5811) );
  CMX2X1 U21666 ( .A0(N7611), .A1(N7610), .S(n3866), .Z(n11523) );
  CMXI2X1 U21667 ( .A0(n11523), .A1(n11517), .S(n4096), .Z(n11530) );
  CMX2X1 U21668 ( .A0(n11518), .A1(n11530), .S(n3812), .Z(n11546) );
  CMXI2X1 U21669 ( .A0(n11519), .A1(n11546), .S(n3432), .Z(N5812) );
  CMX2X1 U21670 ( .A0(N7610), .A1(N7609), .S(n3867), .Z(n11526) );
  CMXI2X1 U21671 ( .A0(n11526), .A1(n11520), .S(n4096), .Z(n11533) );
  CMX2X1 U21672 ( .A0(n11521), .A1(n11533), .S(n4310), .Z(n11549) );
  CMXI2X1 U21673 ( .A0(n11522), .A1(n11549), .S(n3432), .Z(N5813) );
  CMX2X1 U21674 ( .A0(N7609), .A1(N7608), .S(n3864), .Z(n11529) );
  CMXI2X1 U21675 ( .A0(n11529), .A1(n11523), .S(n4096), .Z(n11539) );
  CMX2X1 U21676 ( .A0(n11524), .A1(n11539), .S(n3771), .Z(n11552) );
  CMXI2X1 U21677 ( .A0(n11525), .A1(n11552), .S(n3432), .Z(N5814) );
  CMX2X1 U21678 ( .A0(N7608), .A1(N7607), .S(n3865), .Z(n11532) );
  CMXI2X1 U21679 ( .A0(n11532), .A1(n11526), .S(n4096), .Z(n11542) );
  CMX2X1 U21680 ( .A0(n11527), .A1(n11542), .S(n3772), .Z(n11555) );
  CMXI2X1 U21681 ( .A0(n11528), .A1(n11555), .S(n3432), .Z(N5815) );
  CMX2X1 U21682 ( .A0(N7607), .A1(N7606), .S(n3876), .Z(n11538) );
  CMXI2X1 U21683 ( .A0(n11538), .A1(n11529), .S(n4096), .Z(n11545) );
  CMX2X1 U21684 ( .A0(n11530), .A1(n11545), .S(n3773), .Z(n11558) );
  CMXI2X1 U21685 ( .A0(n11531), .A1(n11558), .S(n3432), .Z(N5816) );
  CMX2X1 U21686 ( .A0(N7606), .A1(N7605), .S(n3877), .Z(n11541) );
  CMXI2X1 U21687 ( .A0(n11541), .A1(n11532), .S(n4096), .Z(n11548) );
  CMX2X1 U21688 ( .A0(n11533), .A1(n11548), .S(n3774), .Z(n11561) );
  CMXI2X1 U21689 ( .A0(n11534), .A1(n11561), .S(n3432), .Z(N5817) );
  CMX2X1 U21690 ( .A0(N8200), .A1(N8199), .S(n3878), .Z(n11601) );
  CMXI2X1 U21691 ( .A0(n11601), .A1(n11535), .S(n4096), .Z(n11668) );
  CMX2X1 U21692 ( .A0(n11536), .A1(n11668), .S(n3775), .Z(n11805) );
  CMXI2X1 U21693 ( .A0(n11537), .A1(n11805), .S(n3432), .Z(N5223) );
  CMX2X1 U21694 ( .A0(N7605), .A1(N7604), .S(n3879), .Z(n11544) );
  CMXI2X1 U21695 ( .A0(n11544), .A1(n11538), .S(n4096), .Z(n11551) );
  CMX2X1 U21696 ( .A0(n11539), .A1(n11551), .S(n3776), .Z(n11564) );
  CMXI2X1 U21697 ( .A0(n11540), .A1(n11564), .S(n3432), .Z(N5818) );
  CMX2X1 U21698 ( .A0(N7604), .A1(N7603), .S(n3876), .Z(n11547) );
  CMXI2X1 U21699 ( .A0(n11547), .A1(n11541), .S(n4096), .Z(n11554) );
  CMX2X1 U21700 ( .A0(n11542), .A1(n11554), .S(n3777), .Z(n11567) );
  CMXI2X1 U21701 ( .A0(n11543), .A1(n11567), .S(n3432), .Z(N5819) );
  CMX2X1 U21702 ( .A0(N7603), .A1(N7602), .S(n3877), .Z(n11550) );
  CMXI2X1 U21703 ( .A0(n11550), .A1(n11544), .S(n4096), .Z(n11557) );
  CMX2X1 U21704 ( .A0(n11545), .A1(n11557), .S(n3790), .Z(n11573) );
  CMXI2X1 U21705 ( .A0(n11546), .A1(n11573), .S(n3431), .Z(N5820) );
  CMX2X1 U21706 ( .A0(N7602), .A1(N7601), .S(n3878), .Z(n11553) );
  CMXI2X1 U21707 ( .A0(n11553), .A1(n11547), .S(n4096), .Z(n11560) );
  CMX2X1 U21708 ( .A0(n11548), .A1(n11560), .S(n3791), .Z(n11576) );
  CMXI2X1 U21709 ( .A0(n11549), .A1(n11576), .S(n3435), .Z(N5821) );
  CMX2X1 U21710 ( .A0(N7601), .A1(N7600), .S(n3879), .Z(n11556) );
  CMXI2X1 U21711 ( .A0(n11556), .A1(n11550), .S(n4095), .Z(n11563) );
  CMX2X1 U21712 ( .A0(n11551), .A1(n11563), .S(n3774), .Z(n11579) );
  CMXI2X1 U21713 ( .A0(n11552), .A1(n11579), .S(n3435), .Z(N5822) );
  CMX2X1 U21714 ( .A0(N7600), .A1(N7599), .S(n3874), .Z(n11559) );
  CMXI2X1 U21715 ( .A0(n11559), .A1(n11553), .S(n4095), .Z(n11566) );
  CMX2X1 U21716 ( .A0(n11554), .A1(n11566), .S(n3810), .Z(n11582) );
  CMXI2X1 U21717 ( .A0(n11555), .A1(n11582), .S(n3434), .Z(N5823) );
  CMX2X1 U21718 ( .A0(N7599), .A1(N7598), .S(n3866), .Z(n11562) );
  CMXI2X1 U21719 ( .A0(n11562), .A1(n11556), .S(n4095), .Z(n11572) );
  CMX2X1 U21720 ( .A0(n11557), .A1(n11572), .S(n3771), .Z(n11585) );
  CMXI2X1 U21721 ( .A0(n11558), .A1(n11585), .S(n3434), .Z(N5824) );
  CMX2X1 U21722 ( .A0(N7598), .A1(N7597), .S(n3867), .Z(n11565) );
  CMXI2X1 U21723 ( .A0(n11565), .A1(n11559), .S(n4095), .Z(n11575) );
  CMX2X1 U21724 ( .A0(n11560), .A1(n11575), .S(n3772), .Z(n11588) );
  CMX2X1 U21725 ( .A0(N7597), .A1(N7596), .S(n3868), .Z(n11571) );
  CMXI2X1 U21726 ( .A0(n11571), .A1(n11562), .S(n4095), .Z(n11578) );
  CMX2X1 U21727 ( .A0(n11563), .A1(n11578), .S(n3773), .Z(n11591) );
  CMX2X1 U21728 ( .A0(N7596), .A1(N7595), .S(n3869), .Z(n11574) );
  CMXI2X1 U21729 ( .A0(n11574), .A1(n11565), .S(n4095), .Z(n11581) );
  CMX2X1 U21730 ( .A0(n11566), .A1(n11581), .S(n3774), .Z(n11594) );
  CMX2X1 U21731 ( .A0(N8199), .A1(N8198), .S(n3870), .Z(n11634) );
  CMXI2X1 U21732 ( .A0(n11634), .A1(n11568), .S(n4095), .Z(n11705) );
  CMX2X1 U21733 ( .A0(n11569), .A1(n11705), .S(n3775), .Z(n11838) );
  CMXI2X1 U21734 ( .A0(n11570), .A1(n11838), .S(n3434), .Z(N5224) );
  CMX2X1 U21735 ( .A0(N7595), .A1(N7594), .S(n3871), .Z(n11577) );
  CMXI2X1 U21736 ( .A0(n11577), .A1(n11571), .S(n4095), .Z(n11584) );
  CMX2X1 U21737 ( .A0(n11572), .A1(n11584), .S(n3810), .Z(n11597) );
  CMX2X1 U21738 ( .A0(N7594), .A1(N7593), .S(n3872), .Z(n11580) );
  CMXI2X1 U21739 ( .A0(n11580), .A1(n11574), .S(n4095), .Z(n11587) );
  CMX2X1 U21740 ( .A0(n11575), .A1(n11587), .S(n3792), .Z(n11600) );
  CMX2X1 U21741 ( .A0(N7593), .A1(N7592), .S(n3868), .Z(n11583) );
  CMXI2X1 U21742 ( .A0(n11583), .A1(n11577), .S(n4095), .Z(n11590) );
  CMX2X1 U21743 ( .A0(n11578), .A1(n11590), .S(n3793), .Z(n11606) );
  CMX2X1 U21744 ( .A0(N7592), .A1(N7591), .S(n3869), .Z(n11586) );
  CMXI2X1 U21745 ( .A0(n11586), .A1(n11580), .S(n4095), .Z(n11593) );
  CMX2X1 U21746 ( .A0(n11581), .A1(n11593), .S(n3794), .Z(n11609) );
  CMX2X1 U21747 ( .A0(N7591), .A1(N7590), .S(n3873), .Z(n11589) );
  CMXI2X1 U21748 ( .A0(n11589), .A1(n11583), .S(n4095), .Z(n11596) );
  CMX2X1 U21749 ( .A0(n11584), .A1(n11596), .S(n3792), .Z(n11612) );
  CMX2X1 U21750 ( .A0(N7590), .A1(N7589), .S(n3874), .Z(n11592) );
  CMXI2X1 U21751 ( .A0(n11592), .A1(n11586), .S(n4095), .Z(n11599) );
  CMX2X1 U21752 ( .A0(n11587), .A1(n11599), .S(n3793), .Z(n11615) );
  CMXI2X1 U21753 ( .A0(n11588), .A1(n11615), .S(n3433), .Z(N5833) );
  CMX2X1 U21754 ( .A0(N7589), .A1(N7588), .S(n3880), .Z(n11595) );
  CMXI2X1 U21755 ( .A0(n11595), .A1(n11589), .S(n4095), .Z(n11605) );
  CMX2X1 U21756 ( .A0(n11590), .A1(n11605), .S(n3794), .Z(n11618) );
  CMXI2X1 U21757 ( .A0(n11591), .A1(n11618), .S(n3433), .Z(N5834) );
  CMX2X1 U21758 ( .A0(N7588), .A1(N7587), .S(n3881), .Z(n11598) );
  CMXI2X1 U21759 ( .A0(n11598), .A1(n11592), .S(n4095), .Z(n11608) );
  CMX2X1 U21760 ( .A0(n11593), .A1(n11608), .S(n3795), .Z(n11621) );
  CMXI2X1 U21761 ( .A0(n11594), .A1(n11621), .S(n3433), .Z(N5835) );
  CMX2X1 U21762 ( .A0(N7587), .A1(N7586), .S(n3862), .Z(n11604) );
  CMXI2X1 U21763 ( .A0(n11604), .A1(n11595), .S(n4095), .Z(n11611) );
  CMX2X1 U21764 ( .A0(n11596), .A1(n11611), .S(n3796), .Z(n11624) );
  CMXI2X1 U21765 ( .A0(n11597), .A1(n11624), .S(n3433), .Z(N5836) );
  CMX2X1 U21766 ( .A0(N7586), .A1(N7585), .S(n3863), .Z(n11607) );
  CMXI2X1 U21767 ( .A0(n11607), .A1(n11598), .S(n4094), .Z(n11614) );
  CMX2X1 U21768 ( .A0(n11599), .A1(n11614), .S(n3797), .Z(n11627) );
  CMXI2X1 U21769 ( .A0(n11600), .A1(n11627), .S(n3433), .Z(N5837) );
  CMX2X1 U21770 ( .A0(N8198), .A1(N8197), .S(n3880), .Z(n11667) );
  CMXI2X1 U21771 ( .A0(n11667), .A1(n11601), .S(n4094), .Z(n11738) );
  CMX2X1 U21772 ( .A0(n11602), .A1(n11738), .S(n3805), .Z(n11871) );
  CMXI2X1 U21773 ( .A0(n11603), .A1(n11871), .S(n3436), .Z(N5225) );
  CMX2X1 U21774 ( .A0(N7585), .A1(N7584), .S(n3881), .Z(n11610) );
  CMXI2X1 U21775 ( .A0(n11610), .A1(n11604), .S(n4094), .Z(n11617) );
  CMX2X1 U21776 ( .A0(n11605), .A1(n11617), .S(n3806), .Z(n11630) );
  CMXI2X1 U21777 ( .A0(n11606), .A1(n11630), .S(n3436), .Z(N5838) );
  CMX2X1 U21778 ( .A0(N7584), .A1(N7583), .S(n3862), .Z(n11613) );
  CMXI2X1 U21779 ( .A0(n11613), .A1(n11607), .S(n4094), .Z(n11620) );
  CMX2X1 U21780 ( .A0(n11608), .A1(n11620), .S(n3807), .Z(n11633) );
  CMXI2X1 U21781 ( .A0(n11609), .A1(n11633), .S(n3436), .Z(N5839) );
  CMX2X1 U21782 ( .A0(N7583), .A1(N7582), .S(n3863), .Z(n11616) );
  CMXI2X1 U21783 ( .A0(n11616), .A1(n11610), .S(n4094), .Z(n11623) );
  CMX2X1 U21784 ( .A0(n11611), .A1(n11623), .S(n3808), .Z(n11639) );
  CMXI2X1 U21785 ( .A0(n11612), .A1(n11639), .S(n3436), .Z(N5840) );
  CMX2X1 U21786 ( .A0(N7582), .A1(N7581), .S(n3875), .Z(n11619) );
  CMXI2X1 U21787 ( .A0(n11619), .A1(n11613), .S(n4094), .Z(n11626) );
  CMX2X1 U21788 ( .A0(n11614), .A1(n11626), .S(n3809), .Z(n11642) );
  CMXI2X1 U21789 ( .A0(n11615), .A1(n11642), .S(n3436), .Z(N5841) );
  CMX2X1 U21790 ( .A0(N7581), .A1(N7580), .S(n3875), .Z(n11622) );
  CMXI2X1 U21791 ( .A0(n11622), .A1(n11616), .S(n4094), .Z(n11629) );
  CMX2X1 U21792 ( .A0(n11617), .A1(n11629), .S(n3810), .Z(n11645) );
  CMXI2X1 U21793 ( .A0(n11618), .A1(n11645), .S(n3436), .Z(N5842) );
  CMX2X1 U21794 ( .A0(N7580), .A1(N7579), .S(n3876), .Z(n11625) );
  CMXI2X1 U21795 ( .A0(n11625), .A1(n11619), .S(n4094), .Z(n11632) );
  CMX2X1 U21796 ( .A0(n11620), .A1(n11632), .S(n3811), .Z(n11648) );
  CMXI2X1 U21797 ( .A0(n11621), .A1(n11648), .S(n3436), .Z(N5843) );
  CMX2X1 U21798 ( .A0(N7579), .A1(N7578), .S(n3877), .Z(n11628) );
  CMXI2X1 U21799 ( .A0(n11628), .A1(n11622), .S(n4094), .Z(n11638) );
  CMX2X1 U21800 ( .A0(n11623), .A1(n11638), .S(n3812), .Z(n11651) );
  CMXI2X1 U21801 ( .A0(n11624), .A1(n11651), .S(n3436), .Z(N5844) );
  CMX2X1 U21802 ( .A0(N7578), .A1(N7577), .S(n3867), .Z(n11631) );
  CMXI2X1 U21803 ( .A0(n11631), .A1(n11625), .S(n4094), .Z(n11641) );
  CMX2X1 U21804 ( .A0(n11626), .A1(n11641), .S(n4363), .Z(n11654) );
  CMXI2X1 U21805 ( .A0(n11627), .A1(n11654), .S(n3436), .Z(N5845) );
  CMX2X1 U21806 ( .A0(N7577), .A1(N7576), .S(n3879), .Z(n11637) );
  CMXI2X1 U21807 ( .A0(n11637), .A1(n11628), .S(n4094), .Z(n11644) );
  CMX2X1 U21808 ( .A0(n11629), .A1(n11644), .S(n3771), .Z(n11657) );
  CMXI2X1 U21809 ( .A0(n11630), .A1(n11657), .S(n3435), .Z(N5846) );
  CMX2X1 U21810 ( .A0(N7576), .A1(N7575), .S(n3880), .Z(n11640) );
  CMXI2X1 U21811 ( .A0(n11640), .A1(n11631), .S(n4094), .Z(n11647) );
  CMX2X1 U21812 ( .A0(n11632), .A1(n11647), .S(n3774), .Z(n11660) );
  CMXI2X1 U21813 ( .A0(n11633), .A1(n11660), .S(n3435), .Z(N5847) );
  CMX2X1 U21814 ( .A0(N8197), .A1(N8196), .S(n3881), .Z(n11704) );
  CMXI2X1 U21815 ( .A0(n11704), .A1(n11634), .S(n4094), .Z(n11771) );
  CMX2X1 U21816 ( .A0(n11635), .A1(n11771), .S(n3775), .Z(n11904) );
  CMXI2X1 U21817 ( .A0(n11636), .A1(n11904), .S(n3435), .Z(N5226) );
  CMX2X1 U21818 ( .A0(N7575), .A1(N7574), .S(n3862), .Z(n11643) );
  CMXI2X1 U21819 ( .A0(n11643), .A1(n11637), .S(n4094), .Z(n11650) );
  CMX2X1 U21820 ( .A0(n11638), .A1(n11650), .S(n3777), .Z(n11663) );
  CMXI2X1 U21821 ( .A0(n11639), .A1(n11663), .S(n3435), .Z(N5848) );
  CMX2X1 U21822 ( .A0(N7574), .A1(N7573), .S(n3863), .Z(n11646) );
  CMXI2X1 U21823 ( .A0(n11646), .A1(n11640), .S(n4094), .Z(n11653) );
  CMX2X1 U21824 ( .A0(n11641), .A1(n11653), .S(n3790), .Z(n11666) );
  CMXI2X1 U21825 ( .A0(n11642), .A1(n11666), .S(n3435), .Z(N5849) );
  CMX2X1 U21826 ( .A0(N7573), .A1(N7572), .S(n3878), .Z(n11649) );
  CMXI2X1 U21827 ( .A0(n11649), .A1(n11643), .S(n4094), .Z(n11656) );
  CMX2X1 U21828 ( .A0(n11644), .A1(n11656), .S(n3791), .Z(n11676) );
  CMXI2X1 U21829 ( .A0(n11645), .A1(n11676), .S(n3435), .Z(N5850) );
  CMX2X1 U21830 ( .A0(N7572), .A1(N7571), .S(n3879), .Z(n11652) );
  CMXI2X1 U21831 ( .A0(n11652), .A1(n11646), .S(n4093), .Z(n11659) );
  CMX2X1 U21832 ( .A0(n11647), .A1(n11659), .S(n3792), .Z(n11679) );
  CMXI2X1 U21833 ( .A0(n11648), .A1(n11679), .S(n3435), .Z(N5851) );
  CMX2X1 U21834 ( .A0(N7571), .A1(N7570), .S(n3868), .Z(n11655) );
  CMXI2X1 U21835 ( .A0(n11655), .A1(n11649), .S(n4093), .Z(n11662) );
  CMX2X1 U21836 ( .A0(n11650), .A1(n11662), .S(n3793), .Z(n11682) );
  CMXI2X1 U21837 ( .A0(n11651), .A1(n11682), .S(n3435), .Z(N5852) );
  CMX2X1 U21838 ( .A0(N7570), .A1(N7569), .S(n3869), .Z(n11658) );
  CMXI2X1 U21839 ( .A0(n11658), .A1(n11652), .S(n4093), .Z(n11665) );
  CMX2X1 U21840 ( .A0(n11653), .A1(n11665), .S(n3807), .Z(n11685) );
  CMXI2X1 U21841 ( .A0(n11654), .A1(n11685), .S(n3435), .Z(N5853) );
  CMX2X1 U21842 ( .A0(N7569), .A1(N7568), .S(n3878), .Z(n11661) );
  CMXI2X1 U21843 ( .A0(n11661), .A1(n11655), .S(n4093), .Z(n11675) );
  CMX2X1 U21844 ( .A0(n11656), .A1(n11675), .S(n3772), .Z(n11688) );
  CMXI2X1 U21845 ( .A0(n11657), .A1(n11688), .S(n3286), .Z(N5854) );
  CMX2X1 U21846 ( .A0(N7568), .A1(N7567), .S(n3879), .Z(n11664) );
  CMXI2X1 U21847 ( .A0(n11664), .A1(n11658), .S(n4093), .Z(n11678) );
  CMX2X1 U21848 ( .A0(n11659), .A1(n11678), .S(n3773), .Z(n11691) );
  CMXI2X1 U21849 ( .A0(n11660), .A1(n11691), .S(n3286), .Z(N5855) );
  CMX2X1 U21850 ( .A0(N7567), .A1(N7566), .S(n3880), .Z(n11674) );
  CMXI2X1 U21851 ( .A0(n11674), .A1(n11661), .S(n4093), .Z(n11681) );
  CMX2X1 U21852 ( .A0(n11662), .A1(n11681), .S(n3806), .Z(n11694) );
  CMXI2X1 U21853 ( .A0(n11663), .A1(n11694), .S(n3286), .Z(N5856) );
  CMX2X1 U21854 ( .A0(N7566), .A1(N7565), .S(n3881), .Z(n11677) );
  CMXI2X1 U21855 ( .A0(n11677), .A1(n11664), .S(n4093), .Z(n11684) );
  CMX2X1 U21856 ( .A0(n11665), .A1(n11684), .S(n3791), .Z(n11697) );
  CMXI2X1 U21857 ( .A0(n11666), .A1(n11697), .S(n3286), .Z(N5857) );
  CMX2X1 U21858 ( .A0(N8196), .A1(N8195), .S(n3862), .Z(n11737) );
  CMXI2X1 U21859 ( .A0(n11737), .A1(n11667), .S(n4093), .Z(n11804) );
  CMX2X1 U21860 ( .A0(n11668), .A1(n11804), .S(n3792), .Z(n11937) );
  CMXI2X1 U21861 ( .A0(n11669), .A1(n11937), .S(n3286), .Z(N5227) );
  CMXI2X1 U21862 ( .A0(n4421), .A1(n11671), .S(n3784), .Z(n11673) );
  CMXI2X1 U21863 ( .A0(n11673), .A1(n11672), .S(n3286), .Z(N5164) );
  CMX2X1 U21864 ( .A0(N7565), .A1(N7564), .S(n3863), .Z(n11680) );
  CMXI2X1 U21865 ( .A0(n11680), .A1(n11674), .S(n4093), .Z(n11687) );
  CMX2X1 U21866 ( .A0(n11675), .A1(n11687), .S(n3793), .Z(n11700) );
  CMXI2X1 U21867 ( .A0(n11676), .A1(n11700), .S(n3286), .Z(N5858) );
  CMXI2X1 U21868 ( .A0(n11683), .A1(n11677), .S(n4093), .Z(n11690) );
  CMX2X1 U21869 ( .A0(n11678), .A1(n11690), .S(n3794), .Z(n11703) );
  CMXI2X1 U21870 ( .A0(n11679), .A1(n11703), .S(n3286), .Z(N5859) );
  CMX2X1 U21871 ( .A0(N7563), .A1(N7562), .S(n3865), .Z(n11686) );
  CMXI2X1 U21872 ( .A0(n11686), .A1(n11680), .S(n4093), .Z(n11693) );
  CMX2X1 U21873 ( .A0(n11681), .A1(n11693), .S(n3795), .Z(n11709) );
  CMXI2X1 U21874 ( .A0(n11682), .A1(n11709), .S(n3286), .Z(N5860) );
  CMX2X1 U21875 ( .A0(N7562), .A1(N7561), .S(n3878), .Z(n11689) );
  CMXI2X1 U21876 ( .A0(n11689), .A1(n11683), .S(n4093), .Z(n11696) );
  CMX2X1 U21877 ( .A0(n11684), .A1(n11696), .S(n3774), .Z(n11712) );
  CMXI2X1 U21878 ( .A0(n11685), .A1(n11712), .S(n3286), .Z(N5861) );
  CMX2X1 U21879 ( .A0(N7561), .A1(N7560), .S(n3870), .Z(n11692) );
  CMXI2X1 U21880 ( .A0(n11692), .A1(n11686), .S(n4093), .Z(n11699) );
  CMX2X1 U21881 ( .A0(n11687), .A1(n11699), .S(n3807), .Z(n11715) );
  CMXI2X1 U21882 ( .A0(n11688), .A1(n11715), .S(n3286), .Z(N5862) );
  CMX2X1 U21883 ( .A0(N7560), .A1(N7559), .S(n3871), .Z(n11695) );
  CMXI2X1 U21884 ( .A0(n11695), .A1(n11689), .S(n4093), .Z(n11702) );
  CMX2X1 U21885 ( .A0(n11690), .A1(n11702), .S(n3808), .Z(n11718) );
  CMXI2X1 U21886 ( .A0(n11691), .A1(n11718), .S(n3411), .Z(N5863) );
  CMX2X1 U21887 ( .A0(N7559), .A1(N7558), .S(n3872), .Z(n11698) );
  CMXI2X1 U21888 ( .A0(n11698), .A1(n11692), .S(n4093), .Z(n11708) );
  CMX2X1 U21889 ( .A0(n11693), .A1(n11708), .S(n3809), .Z(n11721) );
  CMXI2X1 U21890 ( .A0(n11694), .A1(n11721), .S(n3462), .Z(N5864) );
  CMX2X1 U21891 ( .A0(N7558), .A1(N7557), .S(n3873), .Z(n11701) );
  CMXI2X1 U21892 ( .A0(n11701), .A1(n11695), .S(n4093), .Z(n11711) );
  CMX2X1 U21893 ( .A0(n11696), .A1(n11711), .S(n3810), .Z(n11724) );
  CMXI2X1 U21894 ( .A0(n11697), .A1(n11724), .S(n3460), .Z(N5865) );
  CMX2X1 U21895 ( .A0(N7557), .A1(N7556), .S(n3874), .Z(n11707) );
  CMXI2X1 U21896 ( .A0(n11707), .A1(n11698), .S(n4092), .Z(n11714) );
  CMX2X1 U21897 ( .A0(n11699), .A1(n11714), .S(n3811), .Z(n11727) );
  CMXI2X1 U21898 ( .A0(n11700), .A1(n11727), .S(n3459), .Z(N5866) );
  CMX2X1 U21899 ( .A0(N7556), .A1(N7555), .S(n3875), .Z(n11710) );
  CMXI2X1 U21900 ( .A0(n11710), .A1(n11701), .S(n4092), .Z(n11717) );
  CMX2X1 U21901 ( .A0(n11702), .A1(n11717), .S(n3812), .Z(n11730) );
  CMXI2X1 U21902 ( .A0(n11703), .A1(n11730), .S(n3458), .Z(N5867) );
  CMX2X1 U21903 ( .A0(N8195), .A1(N8194), .S(n3876), .Z(n11770) );
  CMXI2X1 U21904 ( .A0(n11770), .A1(n11704), .S(n4092), .Z(n11837) );
  CMX2X1 U21905 ( .A0(n11705), .A1(n11837), .S(n4314), .Z(n11970) );
  CMXI2X1 U21906 ( .A0(n11706), .A1(n11970), .S(n3452), .Z(N5228) );
  CMX2X1 U21907 ( .A0(N7555), .A1(N7554), .S(n3880), .Z(n11713) );
  CMXI2X1 U21908 ( .A0(n11713), .A1(n11707), .S(n4092), .Z(n11720) );
  CMX2X1 U21909 ( .A0(n11708), .A1(n11720), .S(n3771), .Z(n11733) );
  CMXI2X1 U21910 ( .A0(n11709), .A1(n11733), .S(n3457), .Z(N5868) );
  CMX2X1 U21911 ( .A0(N7554), .A1(N7553), .S(n3881), .Z(n11716) );
  CMXI2X1 U21912 ( .A0(n11716), .A1(n11710), .S(n4092), .Z(n11723) );
  CMX2X1 U21913 ( .A0(n11711), .A1(n11723), .S(n3772), .Z(n11736) );
  CMXI2X1 U21914 ( .A0(n11712), .A1(n11736), .S(n3456), .Z(N5869) );
  CMX2X1 U21915 ( .A0(N7553), .A1(N7552), .S(n3880), .Z(n11719) );
  CMXI2X1 U21916 ( .A0(n11719), .A1(n11713), .S(n4092), .Z(n11726) );
  CMX2X1 U21917 ( .A0(n11714), .A1(n11726), .S(n3773), .Z(n11742) );
  CMXI2X1 U21918 ( .A0(n11715), .A1(n11742), .S(n3454), .Z(N5870) );
  CMX2X1 U21919 ( .A0(N7552), .A1(N7551), .S(n3881), .Z(n11722) );
  CMXI2X1 U21920 ( .A0(n11722), .A1(n11716), .S(n4092), .Z(n11729) );
  CMX2X1 U21921 ( .A0(n11717), .A1(n11729), .S(n3774), .Z(n11745) );
  CMXI2X1 U21922 ( .A0(n11718), .A1(n11745), .S(n3453), .Z(N5871) );
  CMX2X1 U21923 ( .A0(N7551), .A1(N7550), .S(n3862), .Z(n11725) );
  CMXI2X1 U21924 ( .A0(n11725), .A1(n11719), .S(n4092), .Z(n11732) );
  CMX2X1 U21925 ( .A0(n11720), .A1(n11732), .S(n3775), .Z(n11748) );
  CMXI2X1 U21926 ( .A0(n11721), .A1(n11748), .S(n3440), .Z(N5872) );
  CMX2X1 U21927 ( .A0(N7550), .A1(N7549), .S(n3863), .Z(n11728) );
  CMXI2X1 U21928 ( .A0(n11728), .A1(n11722), .S(n4092), .Z(n11735) );
  CMX2X1 U21929 ( .A0(n11723), .A1(n11735), .S(n3776), .Z(n11751) );
  CMXI2X1 U21930 ( .A0(n11724), .A1(n11751), .S(n3438), .Z(N5873) );
  CMX2X1 U21931 ( .A0(N7549), .A1(N7548), .S(n3880), .Z(n11731) );
  CMXI2X1 U21932 ( .A0(n11731), .A1(n11725), .S(n4092), .Z(n11741) );
  CMX2X1 U21933 ( .A0(n11726), .A1(n11741), .S(n3777), .Z(n11754) );
  CMXI2X1 U21934 ( .A0(n11727), .A1(n11754), .S(n3437), .Z(N5874) );
  CMX2X1 U21935 ( .A0(N7548), .A1(N7547), .S(n3880), .Z(n11734) );
  CMXI2X1 U21936 ( .A0(n11734), .A1(n11728), .S(n4092), .Z(n11744) );
  CMX2X1 U21937 ( .A0(n11729), .A1(n11744), .S(n3790), .Z(n11757) );
  CMXI2X1 U21938 ( .A0(n11730), .A1(n11757), .S(n3405), .Z(N5875) );
  CMX2X1 U21939 ( .A0(N7547), .A1(N7546), .S(n3881), .Z(n11740) );
  CMXI2X1 U21940 ( .A0(n11740), .A1(n11731), .S(n4092), .Z(n11747) );
  CMX2X1 U21941 ( .A0(n11732), .A1(n11747), .S(n3791), .Z(n11760) );
  CMXI2X1 U21942 ( .A0(n11733), .A1(n11760), .S(n3405), .Z(N5876) );
  CMX2X1 U21943 ( .A0(N7546), .A1(N7545), .S(n3862), .Z(n11743) );
  CMXI2X1 U21944 ( .A0(n11743), .A1(n11734), .S(n4092), .Z(n11750) );
  CMX2X1 U21945 ( .A0(n11735), .A1(n11750), .S(n3797), .Z(n11763) );
  CMXI2X1 U21946 ( .A0(n11736), .A1(n11763), .S(n3405), .Z(N5877) );
  CMX2X1 U21947 ( .A0(N8194), .A1(N8193), .S(n3863), .Z(n11803) );
  CMXI2X1 U21948 ( .A0(n11803), .A1(n11737), .S(n4092), .Z(n11870) );
  CMX2X1 U21949 ( .A0(n11738), .A1(n11870), .S(n3805), .Z(n12003) );
  CMXI2X1 U21950 ( .A0(n11739), .A1(n12003), .S(n3405), .Z(N5229) );
  CMX2X1 U21951 ( .A0(N7545), .A1(N7544), .S(n3864), .Z(n11746) );
  CMXI2X1 U21952 ( .A0(n11746), .A1(n11740), .S(n4092), .Z(n11753) );
  CMX2X1 U21953 ( .A0(n11741), .A1(n11753), .S(n3796), .Z(n11766) );
  CMXI2X1 U21954 ( .A0(n11742), .A1(n11766), .S(n3405), .Z(N5878) );
  CMX2X1 U21955 ( .A0(N7544), .A1(N7543), .S(n3865), .Z(n11749) );
  CMXI2X1 U21956 ( .A0(n11749), .A1(n11743), .S(n4092), .Z(n11756) );
  CMX2X1 U21957 ( .A0(n11744), .A1(n11756), .S(n3797), .Z(n11769) );
  CMXI2X1 U21958 ( .A0(n11745), .A1(n11769), .S(n3405), .Z(N5879) );
  CMX2X1 U21959 ( .A0(N7543), .A1(N7542), .S(n3866), .Z(n11752) );
  CMXI2X1 U21960 ( .A0(n11752), .A1(n11746), .S(n4091), .Z(n11759) );
  CMX2X1 U21961 ( .A0(n11747), .A1(n11759), .S(n3805), .Z(n11775) );
  CMXI2X1 U21962 ( .A0(n11748), .A1(n11775), .S(n3405), .Z(N5880) );
  CMX2X1 U21963 ( .A0(N7542), .A1(N7541), .S(n3880), .Z(n11755) );
  CMXI2X1 U21964 ( .A0(n11755), .A1(n11749), .S(n4091), .Z(n11762) );
  CMX2X1 U21965 ( .A0(n11750), .A1(n11762), .S(n3806), .Z(n11778) );
  CMXI2X1 U21966 ( .A0(n11751), .A1(n11778), .S(n3405), .Z(N5881) );
  CMX2X1 U21967 ( .A0(N7541), .A1(N7540), .S(n3881), .Z(n11758) );
  CMXI2X1 U21968 ( .A0(n11758), .A1(n11752), .S(n4091), .Z(n11765) );
  CMX2X1 U21969 ( .A0(n11753), .A1(n11765), .S(n3807), .Z(n11781) );
  CMXI2X1 U21970 ( .A0(n11754), .A1(n11781), .S(n3404), .Z(N5882) );
  CMX2X1 U21971 ( .A0(N7540), .A1(N7539), .S(n3867), .Z(n11761) );
  CMXI2X1 U21972 ( .A0(n11761), .A1(n11755), .S(n4091), .Z(n11768) );
  CMX2X1 U21973 ( .A0(n11756), .A1(n11768), .S(n3775), .Z(n11784) );
  CMXI2X1 U21974 ( .A0(n11757), .A1(n11784), .S(n3404), .Z(N5883) );
  CMX2X1 U21975 ( .A0(N7539), .A1(N7538), .S(n3868), .Z(n11764) );
  CMXI2X1 U21976 ( .A0(n11764), .A1(n11758), .S(n4091), .Z(n11774) );
  CMX2X1 U21977 ( .A0(n11759), .A1(n11774), .S(n3792), .Z(n11787) );
  CMXI2X1 U21978 ( .A0(n11760), .A1(n11787), .S(n3404), .Z(N5884) );
  CMX2X1 U21979 ( .A0(N7538), .A1(N7537), .S(n3864), .Z(n11767) );
  CMXI2X1 U21980 ( .A0(n11767), .A1(n11761), .S(n4091), .Z(n11777) );
  CMX2X1 U21981 ( .A0(n11762), .A1(n11777), .S(n3793), .Z(n11790) );
  CMXI2X1 U21982 ( .A0(n11763), .A1(n11790), .S(n3404), .Z(N5885) );
  CMX2X1 U21983 ( .A0(N7537), .A1(N7536), .S(n3865), .Z(n11773) );
  CMXI2X1 U21984 ( .A0(n11773), .A1(n11764), .S(n4091), .Z(n11780) );
  CMX2X1 U21985 ( .A0(n11765), .A1(n11780), .S(n3794), .Z(n11793) );
  CMXI2X1 U21986 ( .A0(n11766), .A1(n11793), .S(n3404), .Z(N5886) );
  CMX2X1 U21987 ( .A0(N7536), .A1(N7535), .S(n3866), .Z(n11776) );
  CMXI2X1 U21988 ( .A0(n11776), .A1(n11767), .S(n4091), .Z(n11783) );
  CMX2X1 U21989 ( .A0(n11768), .A1(n11783), .S(n3795), .Z(n11796) );
  CMXI2X1 U21990 ( .A0(n11769), .A1(n11796), .S(n3404), .Z(N5887) );
  CMX2X1 U21991 ( .A0(N8193), .A1(N8192), .S(n3867), .Z(n11836) );
  CMXI2X1 U21992 ( .A0(n11836), .A1(n11770), .S(n4091), .Z(n11903) );
  CMX2X1 U21993 ( .A0(n11771), .A1(n11903), .S(n3796), .Z(n12040) );
  CMXI2X1 U21994 ( .A0(n11772), .A1(n12040), .S(n3404), .Z(N5230) );
  CMX2X1 U21995 ( .A0(N7535), .A1(N7534), .S(n3864), .Z(n11779) );
  CMXI2X1 U21996 ( .A0(n11779), .A1(n11773), .S(n4091), .Z(n11786) );
  CMX2X1 U21997 ( .A0(n11774), .A1(n11786), .S(n3797), .Z(n11799) );
  CMXI2X1 U21998 ( .A0(n11775), .A1(n11799), .S(n3404), .Z(N5888) );
  CMX2X1 U21999 ( .A0(N7534), .A1(N7533), .S(n3865), .Z(n11782) );
  CMXI2X1 U22000 ( .A0(n11782), .A1(n11776), .S(n4091), .Z(n11789) );
  CMX2X1 U22001 ( .A0(n11777), .A1(n11789), .S(n3805), .Z(n11802) );
  CMXI2X1 U22002 ( .A0(n11778), .A1(n11802), .S(n3404), .Z(N5889) );
  CMX2X1 U22003 ( .A0(N7533), .A1(N7532), .S(n3866), .Z(n11785) );
  CMXI2X1 U22004 ( .A0(n11785), .A1(n11779), .S(n4091), .Z(n11792) );
  CMX2X1 U22005 ( .A0(n11780), .A1(n11792), .S(n3806), .Z(n11808) );
  CMXI2X1 U22006 ( .A0(n11781), .A1(n11808), .S(n3404), .Z(N5890) );
  CMX2X1 U22007 ( .A0(N7532), .A1(N7531), .S(n3867), .Z(n11788) );
  CMXI2X1 U22008 ( .A0(n11788), .A1(n11782), .S(n4091), .Z(n11795) );
  CMX2X1 U22009 ( .A0(n11783), .A1(n11795), .S(n3807), .Z(n11811) );
  CMXI2X1 U22010 ( .A0(n11784), .A1(n11811), .S(n3407), .Z(N5891) );
  CMX2X1 U22011 ( .A0(N7531), .A1(N7530), .S(n3881), .Z(n11791) );
  CMXI2X1 U22012 ( .A0(n11791), .A1(n11785), .S(n4091), .Z(n11798) );
  CMX2X1 U22013 ( .A0(n11786), .A1(n11798), .S(n3808), .Z(n11814) );
  CMXI2X1 U22014 ( .A0(n11787), .A1(n11814), .S(n3407), .Z(N5892) );
  CMX2X1 U22015 ( .A0(N7530), .A1(N7529), .S(n3869), .Z(n11794) );
  CMXI2X1 U22016 ( .A0(n11794), .A1(n11788), .S(n4091), .Z(n11801) );
  CMX2X1 U22017 ( .A0(n11789), .A1(n11801), .S(n3809), .Z(n11817) );
  CMXI2X1 U22018 ( .A0(n11790), .A1(n11817), .S(n3407), .Z(N5893) );
  CMX2X1 U22019 ( .A0(N7529), .A1(N7528), .S(n3870), .Z(n11797) );
  CMXI2X1 U22020 ( .A0(n11797), .A1(n11791), .S(n4091), .Z(n11807) );
  CMX2X1 U22021 ( .A0(n11792), .A1(n11807), .S(n3810), .Z(n11820) );
  CMXI2X1 U22022 ( .A0(n11793), .A1(n11820), .S(n3407), .Z(N5894) );
  CMX2X1 U22023 ( .A0(N7528), .A1(N7527), .S(n3871), .Z(n11800) );
  CMXI2X1 U22024 ( .A0(n11800), .A1(n11794), .S(n4090), .Z(n11810) );
  CMX2X1 U22025 ( .A0(n11795), .A1(n11810), .S(n3811), .Z(n11823) );
  CMXI2X1 U22026 ( .A0(n11796), .A1(n11823), .S(n3406), .Z(N5895) );
  CMXI2X1 U22027 ( .A0(n11806), .A1(n11797), .S(n4090), .Z(n11813) );
  CMX2X1 U22028 ( .A0(n11798), .A1(n11813), .S(n3812), .Z(n11826) );
  CMXI2X1 U22029 ( .A0(n11799), .A1(n11826), .S(n3406), .Z(N5896) );
  CMX2X1 U22030 ( .A0(N7526), .A1(N7525), .S(n3873), .Z(n11809) );
  CMXI2X1 U22031 ( .A0(n11809), .A1(n11800), .S(n4090), .Z(n11816) );
  CMX2X1 U22032 ( .A0(n11801), .A1(n11816), .S(n4313), .Z(n11829) );
  CMXI2X1 U22033 ( .A0(n11802), .A1(n11829), .S(n3406), .Z(N5897) );
  CMX2X1 U22034 ( .A0(N8192), .A1(N8191), .S(n3874), .Z(n11869) );
  CMXI2X1 U22035 ( .A0(n11869), .A1(n11803), .S(n4090), .Z(n11936) );
  CMX2X1 U22036 ( .A0(n11804), .A1(n11936), .S(n3773), .Z(n12073) );
  CMXI2X1 U22037 ( .A0(n11805), .A1(n12073), .S(n3406), .Z(N5231) );
  CMX2X1 U22038 ( .A0(N7525), .A1(N7524), .S(n3875), .Z(n11812) );
  CMXI2X1 U22039 ( .A0(n11812), .A1(n11806), .S(n4090), .Z(n11819) );
  CMX2X1 U22040 ( .A0(n11807), .A1(n11819), .S(n3774), .Z(n11832) );
  CMXI2X1 U22041 ( .A0(n11808), .A1(n11832), .S(n3406), .Z(N5898) );
  CMX2X1 U22042 ( .A0(N7524), .A1(N7523), .S(n3862), .Z(n11815) );
  CMXI2X1 U22043 ( .A0(n11815), .A1(n11809), .S(n4090), .Z(n11822) );
  CMX2X1 U22044 ( .A0(n11810), .A1(n11822), .S(n3775), .Z(n11835) );
  CMXI2X1 U22045 ( .A0(n11811), .A1(n11835), .S(n3406), .Z(N5899) );
  CMX2X1 U22046 ( .A0(N7523), .A1(N7522), .S(n3863), .Z(n11818) );
  CMXI2X1 U22047 ( .A0(n11818), .A1(n11812), .S(n4090), .Z(n11825) );
  CMX2X1 U22048 ( .A0(n11813), .A1(n11825), .S(n3776), .Z(n11841) );
  CMXI2X1 U22049 ( .A0(n11814), .A1(n11841), .S(n3406), .Z(N5900) );
  CMX2X1 U22050 ( .A0(N7522), .A1(N7521), .S(n3876), .Z(n11821) );
  CMXI2X1 U22051 ( .A0(n11821), .A1(n11815), .S(n4090), .Z(n11828) );
  CMX2X1 U22052 ( .A0(n11816), .A1(n11828), .S(n3777), .Z(n11844) );
  CMXI2X1 U22053 ( .A0(n11817), .A1(n11844), .S(n3406), .Z(N5901) );
  CMX2X1 U22054 ( .A0(N7521), .A1(N7520), .S(n3877), .Z(n11824) );
  CMXI2X1 U22055 ( .A0(n11824), .A1(n11818), .S(n4090), .Z(n11831) );
  CMX2X1 U22056 ( .A0(n11819), .A1(n11831), .S(n3790), .Z(n11847) );
  CMXI2X1 U22057 ( .A0(n11820), .A1(n11847), .S(n3406), .Z(N5902) );
  CMX2X1 U22058 ( .A0(N7520), .A1(N7519), .S(n3868), .Z(n11827) );
  CMXI2X1 U22059 ( .A0(n11827), .A1(n11821), .S(n4090), .Z(n11834) );
  CMX2X1 U22060 ( .A0(n11822), .A1(n11834), .S(n3791), .Z(n11850) );
  CMXI2X1 U22061 ( .A0(n11823), .A1(n11850), .S(n3406), .Z(N5903) );
  CMX2X1 U22062 ( .A0(N7519), .A1(N7518), .S(n3869), .Z(n11830) );
  CMXI2X1 U22063 ( .A0(n11830), .A1(n11824), .S(n4090), .Z(n11840) );
  CMX2X1 U22064 ( .A0(n11825), .A1(n11840), .S(n3792), .Z(n11853) );
  CMXI2X1 U22065 ( .A0(n11826), .A1(n11853), .S(n3406), .Z(N5904) );
  CMX2X1 U22066 ( .A0(N7518), .A1(N7517), .S(n3870), .Z(n11833) );
  CMXI2X1 U22067 ( .A0(n11833), .A1(n11827), .S(n4090), .Z(n11843) );
  CMX2X1 U22068 ( .A0(n11828), .A1(n11843), .S(n3793), .Z(n11856) );
  CMXI2X1 U22069 ( .A0(n11829), .A1(n11856), .S(n3405), .Z(N5905) );
  CMX2X1 U22070 ( .A0(N7517), .A1(N7516), .S(n3871), .Z(n11839) );
  CMXI2X1 U22071 ( .A0(n11839), .A1(n11830), .S(n4090), .Z(n11846) );
  CMX2X1 U22072 ( .A0(n11831), .A1(n11846), .S(n3794), .Z(n11859) );
  CMXI2X1 U22073 ( .A0(n11832), .A1(n11859), .S(n3405), .Z(N5906) );
  CMX2X1 U22074 ( .A0(N7516), .A1(N7515), .S(n3868), .Z(n11842) );
  CMXI2X1 U22075 ( .A0(n11842), .A1(n11833), .S(n4090), .Z(n11849) );
  CMX2X1 U22076 ( .A0(n11834), .A1(n11849), .S(n3795), .Z(n11862) );
  CMXI2X1 U22077 ( .A0(n11835), .A1(n11862), .S(n3405), .Z(N5907) );
  CMX2X1 U22078 ( .A0(N8191), .A1(N8190), .S(n3869), .Z(n11902) );
  CMXI2X1 U22079 ( .A0(n11902), .A1(n11836), .S(n4090), .Z(n11969) );
  CMX2X1 U22080 ( .A0(n11837), .A1(n11969), .S(n3796), .Z(n12106) );
  CMXI2X1 U22081 ( .A0(n11838), .A1(n12106), .S(n3408), .Z(N5232) );
  CMX2X1 U22082 ( .A0(N7515), .A1(N7514), .S(n3870), .Z(n11845) );
  CMXI2X1 U22083 ( .A0(n11845), .A1(n11839), .S(n4090), .Z(n11852) );
  CMX2X1 U22084 ( .A0(n11840), .A1(n11852), .S(n3797), .Z(n11865) );
  CMXI2X1 U22085 ( .A0(n11841), .A1(n11865), .S(n3408), .Z(N5908) );
  CMX2X1 U22086 ( .A0(N7514), .A1(N7513), .S(n3871), .Z(n11848) );
  CMXI2X1 U22087 ( .A0(n11848), .A1(n11842), .S(n4089), .Z(n11855) );
  CMX2X1 U22088 ( .A0(n11843), .A1(n11855), .S(n3805), .Z(n11868) );
  CMXI2X1 U22089 ( .A0(n11844), .A1(n11868), .S(n3408), .Z(N5909) );
  CMX2X1 U22090 ( .A0(N7513), .A1(N7512), .S(n3862), .Z(n11851) );
  CMXI2X1 U22091 ( .A0(n11851), .A1(n11845), .S(n4089), .Z(n11858) );
  CMX2X1 U22092 ( .A0(n11846), .A1(n11858), .S(n3806), .Z(n11874) );
  CMXI2X1 U22093 ( .A0(n11847), .A1(n11874), .S(n3408), .Z(N5910) );
  CMX2X1 U22094 ( .A0(N7512), .A1(N7511), .S(n3878), .Z(n11854) );
  CMXI2X1 U22095 ( .A0(n11854), .A1(n11848), .S(n4089), .Z(n11861) );
  CMX2X1 U22096 ( .A0(n11849), .A1(n11861), .S(n3776), .Z(n11877) );
  CMXI2X1 U22097 ( .A0(n11850), .A1(n11877), .S(n3408), .Z(N5911) );
  CMX2X1 U22098 ( .A0(N7511), .A1(N7510), .S(n3879), .Z(n11857) );
  CMXI2X1 U22099 ( .A0(n11857), .A1(n11851), .S(n4089), .Z(n11864) );
  CMX2X1 U22100 ( .A0(n11852), .A1(n11864), .S(n3812), .Z(n11880) );
  CMXI2X1 U22101 ( .A0(n11853), .A1(n11880), .S(n3408), .Z(N5912) );
  CMX2X1 U22102 ( .A0(N7510), .A1(N7509), .S(n3880), .Z(n11860) );
  CMXI2X1 U22103 ( .A0(n11860), .A1(n11854), .S(n4089), .Z(n11867) );
  CMX2X1 U22104 ( .A0(n11855), .A1(n11867), .S(n3793), .Z(n11883) );
  CMXI2X1 U22105 ( .A0(n11856), .A1(n11883), .S(n3408), .Z(N5913) );
  CMX2X1 U22106 ( .A0(N7509), .A1(N7508), .S(n3881), .Z(n11863) );
  CMXI2X1 U22107 ( .A0(n11863), .A1(n11857), .S(n4089), .Z(n11873) );
  CMX2X1 U22108 ( .A0(n11858), .A1(n11873), .S(n3794), .Z(n11886) );
  CMXI2X1 U22109 ( .A0(n11859), .A1(n11886), .S(n3408), .Z(N5914) );
  CMX2X1 U22110 ( .A0(N7508), .A1(N7507), .S(n3862), .Z(n11866) );
  CMXI2X1 U22111 ( .A0(n11866), .A1(n11860), .S(n4089), .Z(n11876) );
  CMX2X1 U22112 ( .A0(n11861), .A1(n11876), .S(n3795), .Z(n11889) );
  CMXI2X1 U22113 ( .A0(n11862), .A1(n11889), .S(n3408), .Z(N5915) );
  CMX2X1 U22114 ( .A0(N7507), .A1(N7506), .S(n3863), .Z(n11872) );
  CMXI2X1 U22115 ( .A0(n11872), .A1(n11863), .S(n4089), .Z(n11879) );
  CMX2X1 U22116 ( .A0(n11864), .A1(n11879), .S(n3796), .Z(n11892) );
  CMXI2X1 U22117 ( .A0(n11865), .A1(n11892), .S(n3408), .Z(N5916) );
  CMX2X1 U22118 ( .A0(N7506), .A1(N7505), .S(n3864), .Z(n11875) );
  CMXI2X1 U22119 ( .A0(n11875), .A1(n11866), .S(n4089), .Z(n11882) );
  CMX2X1 U22120 ( .A0(n11867), .A1(n11882), .S(n3797), .Z(n11895) );
  CMXI2X1 U22121 ( .A0(n11868), .A1(n11895), .S(n3408), .Z(N5917) );
  CMX2X1 U22122 ( .A0(N8190), .A1(N8189), .S(n3864), .Z(n11935) );
  CMXI2X1 U22123 ( .A0(n11935), .A1(n11869), .S(n4089), .Z(n12002) );
  CMX2X1 U22124 ( .A0(n11870), .A1(n12002), .S(n3795), .Z(n12139) );
  CMXI2X1 U22125 ( .A0(n11871), .A1(n12139), .S(n3407), .Z(N5233) );
  CMX2X1 U22126 ( .A0(N7505), .A1(N7504), .S(n3865), .Z(n11878) );
  CMXI2X1 U22127 ( .A0(n11878), .A1(n11872), .S(n4089), .Z(n11885) );
  CMX2X1 U22128 ( .A0(n11873), .A1(n11885), .S(n3796), .Z(n11898) );
  CMXI2X1 U22129 ( .A0(n11874), .A1(n11898), .S(n3407), .Z(N5918) );
  CMX2X1 U22130 ( .A0(N7504), .A1(N7503), .S(n3865), .Z(n11881) );
  CMXI2X1 U22131 ( .A0(n11881), .A1(n11875), .S(n4089), .Z(n11888) );
  CMX2X1 U22132 ( .A0(n11876), .A1(n11888), .S(n3797), .Z(n11901) );
  CMXI2X1 U22133 ( .A0(n11877), .A1(n11901), .S(n3407), .Z(N5919) );
  CMX2X1 U22134 ( .A0(N7503), .A1(N7502), .S(n3866), .Z(n11884) );
  CMXI2X1 U22135 ( .A0(n11884), .A1(n11878), .S(n4089), .Z(n11891) );
  CMX2X1 U22136 ( .A0(n11879), .A1(n11891), .S(n3805), .Z(n11907) );
  CMXI2X1 U22137 ( .A0(n11880), .A1(n11907), .S(n3407), .Z(N5920) );
  CMX2X1 U22138 ( .A0(N7502), .A1(N7501), .S(n3872), .Z(n11887) );
  CMXI2X1 U22139 ( .A0(n11887), .A1(n11881), .S(n4089), .Z(n11894) );
  CMX2X1 U22140 ( .A0(n11882), .A1(n11894), .S(n3806), .Z(n11910) );
  CMXI2X1 U22141 ( .A0(n11883), .A1(n11910), .S(n3407), .Z(N5921) );
  CMX2X1 U22142 ( .A0(N7501), .A1(N7500), .S(n3873), .Z(n11890) );
  CMXI2X1 U22143 ( .A0(n11890), .A1(n11884), .S(n4089), .Z(n11897) );
  CMX2X1 U22144 ( .A0(n11885), .A1(n11897), .S(n3807), .Z(n11913) );
  CMXI2X1 U22145 ( .A0(n11886), .A1(n11913), .S(n3407), .Z(N5922) );
  CMX2X1 U22146 ( .A0(N7500), .A1(N7499), .S(n3874), .Z(n11893) );
  CMXI2X1 U22147 ( .A0(n11893), .A1(n11887), .S(n4089), .Z(n11900) );
  CMX2X1 U22148 ( .A0(n11888), .A1(n11900), .S(n3808), .Z(n11916) );
  CMXI2X1 U22149 ( .A0(n11889), .A1(n11916), .S(n3407), .Z(N5923) );
  CMX2X1 U22150 ( .A0(N7499), .A1(N7498), .S(n3875), .Z(n11896) );
  CMXI2X1 U22151 ( .A0(n11896), .A1(n11890), .S(n4088), .Z(n11906) );
  CMX2X1 U22152 ( .A0(n11891), .A1(n11906), .S(n3809), .Z(n11919) );
  CMXI2X1 U22153 ( .A0(n11892), .A1(n11919), .S(n3410), .Z(N5924) );
  CMX2X1 U22154 ( .A0(N7498), .A1(N7497), .S(n3872), .Z(n11899) );
  CMXI2X1 U22155 ( .A0(n11899), .A1(n11893), .S(n4088), .Z(n11909) );
  CMX2X1 U22156 ( .A0(n11894), .A1(n11909), .S(n3810), .Z(n11922) );
  CMXI2X1 U22157 ( .A0(n11895), .A1(n11922), .S(n3410), .Z(N5925) );
  CMX2X1 U22158 ( .A0(N7497), .A1(N7496), .S(n3873), .Z(n11905) );
  CMXI2X1 U22159 ( .A0(n11905), .A1(n11896), .S(n4088), .Z(n11912) );
  CMX2X1 U22160 ( .A0(n11897), .A1(n11912), .S(n3811), .Z(n11925) );
  CMXI2X1 U22161 ( .A0(n11898), .A1(n11925), .S(n3410), .Z(N5926) );
  CMX2X1 U22162 ( .A0(N7496), .A1(N7495), .S(n3874), .Z(n11908) );
  CMXI2X1 U22163 ( .A0(n11908), .A1(n11899), .S(n4088), .Z(n11915) );
  CMX2X1 U22164 ( .A0(n11900), .A1(n11915), .S(n3812), .Z(n11928) );
  CMXI2X1 U22165 ( .A0(n11901), .A1(n11928), .S(n3410), .Z(N5927) );
  CMX2X1 U22166 ( .A0(N8189), .A1(N8188), .S(n3875), .Z(n11968) );
  CMXI2X1 U22167 ( .A0(n11968), .A1(n11902), .S(n4088), .Z(n12039) );
  CMX2X1 U22168 ( .A0(n11903), .A1(n12039), .S(n4317), .Z(n12172) );
  CMXI2X1 U22169 ( .A0(n11904), .A1(n12172), .S(n3410), .Z(N5234) );
  CMX2X1 U22170 ( .A0(N7495), .A1(N7494), .S(n3863), .Z(n11911) );
  CMXI2X1 U22171 ( .A0(n11911), .A1(n11905), .S(n4088), .Z(n11918) );
  CMX2X1 U22172 ( .A0(n11906), .A1(n11918), .S(n3771), .Z(n11931) );
  CMXI2X1 U22173 ( .A0(n11907), .A1(n11931), .S(n3410), .Z(N5928) );
  CMX2X1 U22174 ( .A0(N7494), .A1(N7493), .S(n3867), .Z(n11914) );
  CMXI2X1 U22175 ( .A0(n11914), .A1(n11908), .S(n4088), .Z(n11921) );
  CMX2X1 U22176 ( .A0(n11909), .A1(n11921), .S(n3792), .Z(n11934) );
  CMXI2X1 U22177 ( .A0(n11910), .A1(n11934), .S(n3410), .Z(N5929) );
  CMX2X1 U22178 ( .A0(N7493), .A1(N7492), .S(n3868), .Z(n11917) );
  CMXI2X1 U22179 ( .A0(n11917), .A1(n11911), .S(n4088), .Z(n11924) );
  CMX2X1 U22180 ( .A0(n11912), .A1(n11924), .S(n3793), .Z(n11940) );
  CMXI2X1 U22181 ( .A0(n11913), .A1(n11940), .S(n3409), .Z(N5930) );
  CMX2X1 U22182 ( .A0(N7492), .A1(N7491), .S(n3870), .Z(n11920) );
  CMXI2X1 U22183 ( .A0(n11920), .A1(n11914), .S(n4088), .Z(n11927) );
  CMX2X1 U22184 ( .A0(n11915), .A1(n11927), .S(n3795), .Z(n11943) );
  CMXI2X1 U22185 ( .A0(n11916), .A1(n11943), .S(n3409), .Z(N5931) );
  CMX2X1 U22186 ( .A0(N7491), .A1(N7490), .S(n3871), .Z(n11923) );
  CMXI2X1 U22187 ( .A0(n11923), .A1(n11917), .S(n4088), .Z(n11930) );
  CMX2X1 U22188 ( .A0(n11918), .A1(n11930), .S(n3796), .Z(n11946) );
  CMXI2X1 U22189 ( .A0(n11919), .A1(n11946), .S(n3409), .Z(N5932) );
  CMX2X1 U22190 ( .A0(N7490), .A1(N7489), .S(n3872), .Z(n11926) );
  CMXI2X1 U22191 ( .A0(n11926), .A1(n11920), .S(n4088), .Z(n11933) );
  CMX2X1 U22192 ( .A0(n11921), .A1(n11933), .S(n3797), .Z(n11949) );
  CMXI2X1 U22193 ( .A0(n11922), .A1(n11949), .S(n3409), .Z(N5933) );
  CMX2X1 U22194 ( .A0(N7489), .A1(N7488), .S(n3873), .Z(n11929) );
  CMXI2X1 U22195 ( .A0(n11929), .A1(n11923), .S(n4088), .Z(n11939) );
  CMX2X1 U22196 ( .A0(n11924), .A1(n11939), .S(n3805), .Z(n11952) );
  CMXI2X1 U22197 ( .A0(n11925), .A1(n11952), .S(n3409), .Z(N5934) );
  CMX2X1 U22198 ( .A0(N7488), .A1(N7487), .S(n3866), .Z(n11932) );
  CMXI2X1 U22199 ( .A0(n11932), .A1(n11926), .S(n4088), .Z(n11942) );
  CMX2X1 U22200 ( .A0(n11927), .A1(n11942), .S(n3806), .Z(n11955) );
  CMXI2X1 U22201 ( .A0(n11928), .A1(n11955), .S(n3409), .Z(N5935) );
  CMX2X1 U22202 ( .A0(N7487), .A1(N7486), .S(n3867), .Z(n11938) );
  CMXI2X1 U22203 ( .A0(n11938), .A1(n11929), .S(n4088), .Z(n11945) );
  CMX2X1 U22204 ( .A0(n11930), .A1(n11945), .S(n4311), .Z(n11958) );
  CMXI2X1 U22205 ( .A0(n11931), .A1(n11958), .S(n3409), .Z(N5936) );
  CMX2X1 U22206 ( .A0(N7486), .A1(N7485), .S(n3874), .Z(n11941) );
  CMXI2X1 U22207 ( .A0(n11941), .A1(n11932), .S(n4088), .Z(n11948) );
  CMX2X1 U22208 ( .A0(n11933), .A1(n11948), .S(n3772), .Z(n11961) );
  CMXI2X1 U22209 ( .A0(n11934), .A1(n11961), .S(n3409), .Z(N5937) );
  CMX2X1 U22210 ( .A0(N8188), .A1(N8187), .S(n3875), .Z(n12001) );
  CMXI2X1 U22211 ( .A0(n12001), .A1(n11935), .S(n4088), .Z(n12072) );
  CMX2X1 U22212 ( .A0(n11936), .A1(n12072), .S(n3773), .Z(n12205) );
  CMXI2X1 U22213 ( .A0(n11937), .A1(n12205), .S(n3409), .Z(N5235) );
  CMX2X1 U22214 ( .A0(N7485), .A1(N7484), .S(n3876), .Z(n11944) );
  CMXI2X1 U22215 ( .A0(n11944), .A1(n11938), .S(n4087), .Z(n11951) );
  CMX2X1 U22216 ( .A0(n11939), .A1(n11951), .S(n3774), .Z(n11964) );
  CMXI2X1 U22217 ( .A0(n11940), .A1(n11964), .S(n3409), .Z(N5938) );
  CMX2X1 U22218 ( .A0(N7484), .A1(N7483), .S(n3877), .Z(n11947) );
  CMXI2X1 U22219 ( .A0(n11947), .A1(n11941), .S(n4087), .Z(n11954) );
  CMX2X1 U22220 ( .A0(n11942), .A1(n11954), .S(n3775), .Z(n11967) );
  CMXI2X1 U22221 ( .A0(n11943), .A1(n11967), .S(n3409), .Z(N5939) );
  CMX2X1 U22222 ( .A0(N7483), .A1(N7482), .S(n3878), .Z(n11950) );
  CMXI2X1 U22223 ( .A0(n11950), .A1(n11944), .S(n4087), .Z(n11957) );
  CMX2X1 U22224 ( .A0(n11945), .A1(n11957), .S(n3776), .Z(n11973) );
  CMXI2X1 U22225 ( .A0(n11946), .A1(n11973), .S(n3446), .Z(N5940) );
  CMX2X1 U22226 ( .A0(N7482), .A1(N7481), .S(n3879), .Z(n11953) );
  CMXI2X1 U22227 ( .A0(n11953), .A1(n11947), .S(n4087), .Z(n11960) );
  CMX2X1 U22228 ( .A0(n11948), .A1(n11960), .S(n3777), .Z(n11976) );
  CMXI2X1 U22229 ( .A0(n11949), .A1(n11976), .S(n3446), .Z(N5941) );
  CMX2X1 U22230 ( .A0(N7481), .A1(N7480), .S(n3876), .Z(n11956) );
  CMXI2X1 U22231 ( .A0(n11956), .A1(n11950), .S(n4087), .Z(n11963) );
  CMX2X1 U22232 ( .A0(n11951), .A1(n11963), .S(n3791), .Z(n11979) );
  CMXI2X1 U22233 ( .A0(n11952), .A1(n11979), .S(n3455), .Z(N5942) );
  CMX2X1 U22234 ( .A0(N7480), .A1(N7479), .S(n3877), .Z(n11959) );
  CMXI2X1 U22235 ( .A0(n11959), .A1(n11953), .S(n4087), .Z(n11966) );
  CMX2X1 U22236 ( .A0(n11954), .A1(n11966), .S(n3792), .Z(n11982) );
  CMXI2X1 U22237 ( .A0(n11955), .A1(n11982), .S(n3411), .Z(N5943) );
  CMX2X1 U22238 ( .A0(N7479), .A1(N7478), .S(n3878), .Z(n11962) );
  CMXI2X1 U22239 ( .A0(n11962), .A1(n11956), .S(n4087), .Z(n11972) );
  CMX2X1 U22240 ( .A0(n11957), .A1(n11972), .S(n3793), .Z(n11985) );
  CMXI2X1 U22241 ( .A0(n11958), .A1(n11985), .S(n3411), .Z(N5944) );
  CMX2X1 U22242 ( .A0(N7478), .A1(N7477), .S(n3879), .Z(n11965) );
  CMXI2X1 U22243 ( .A0(n11965), .A1(n11959), .S(n4087), .Z(n11975) );
  CMX2X1 U22244 ( .A0(n11960), .A1(n11975), .S(n3794), .Z(n11988) );
  CMXI2X1 U22245 ( .A0(n11961), .A1(n11988), .S(n3411), .Z(N5945) );
  CMX2X1 U22246 ( .A0(N7477), .A1(N7476), .S(n3864), .Z(n11971) );
  CMXI2X1 U22247 ( .A0(n11971), .A1(n11962), .S(n4087), .Z(n11978) );
  CMX2X1 U22248 ( .A0(n11963), .A1(n11978), .S(n3795), .Z(n11991) );
  CMXI2X1 U22249 ( .A0(n11964), .A1(n11991), .S(n3411), .Z(N5946) );
  CMX2X1 U22250 ( .A0(N7476), .A1(N7475), .S(n3876), .Z(n11974) );
  CMXI2X1 U22251 ( .A0(n11974), .A1(n11965), .S(n4087), .Z(n11981) );
  CMX2X1 U22252 ( .A0(n11966), .A1(n11981), .S(n3796), .Z(n11994) );
  CMXI2X1 U22253 ( .A0(n11967), .A1(n11994), .S(n3411), .Z(N5947) );
  CMX2X1 U22254 ( .A0(N8187), .A1(N8186), .S(n3877), .Z(n12038) );
  CMXI2X1 U22255 ( .A0(n12038), .A1(n11968), .S(n4087), .Z(n12105) );
  CMX2X1 U22256 ( .A0(n11969), .A1(n12105), .S(n3797), .Z(n12239) );
  CMXI2X1 U22257 ( .A0(n11970), .A1(n12239), .S(n3411), .Z(N5236) );
  CMX2X1 U22258 ( .A0(N7475), .A1(N7474), .S(n3878), .Z(n11977) );
  CMXI2X1 U22259 ( .A0(n11977), .A1(n11971), .S(n4087), .Z(n11984) );
  CMX2X1 U22260 ( .A0(n11972), .A1(n11984), .S(n3805), .Z(n11997) );
  CMXI2X1 U22261 ( .A0(n11973), .A1(n11997), .S(n3411), .Z(N5948) );
  CMX2X1 U22262 ( .A0(N7474), .A1(N7473), .S(n3879), .Z(n11980) );
  CMXI2X1 U22263 ( .A0(n11980), .A1(n11974), .S(n4087), .Z(n11987) );
  CMX2X1 U22264 ( .A0(n11975), .A1(n11987), .S(n3806), .Z(n12000) );
  CMXI2X1 U22265 ( .A0(n11976), .A1(n12000), .S(n3411), .Z(N5949) );
  CMX2X1 U22266 ( .A0(N7473), .A1(N7472), .S(n3880), .Z(n11983) );
  CMXI2X1 U22267 ( .A0(n11983), .A1(n11977), .S(n4087), .Z(n11990) );
  CMX2X1 U22268 ( .A0(n11978), .A1(n11990), .S(n3793), .Z(n12010) );
  CMXI2X1 U22269 ( .A0(n11979), .A1(n12010), .S(n3411), .Z(N5950) );
  CMX2X1 U22270 ( .A0(N7472), .A1(N7471), .S(n3881), .Z(n11986) );
  CMXI2X1 U22271 ( .A0(n11986), .A1(n11980), .S(n4087), .Z(n11993) );
  CMX2X1 U22272 ( .A0(n11981), .A1(n11993), .S(n3794), .Z(n12013) );
  CMXI2X1 U22273 ( .A0(n11982), .A1(n12013), .S(n3411), .Z(N5951) );
  CMX2X1 U22274 ( .A0(N7471), .A1(N7470), .S(n3862), .Z(n11989) );
  CMXI2X1 U22275 ( .A0(n11989), .A1(n11983), .S(n4087), .Z(n11996) );
  CMX2X1 U22276 ( .A0(n11984), .A1(n11996), .S(n3807), .Z(n12016) );
  CMXI2X1 U22277 ( .A0(n11985), .A1(n12016), .S(n3410), .Z(N5952) );
  CMX2X1 U22278 ( .A0(N7470), .A1(N7469), .S(n3868), .Z(n11992) );
  CMXI2X1 U22279 ( .A0(n11992), .A1(n11986), .S(n4086), .Z(n11999) );
  CMX2X1 U22280 ( .A0(n11987), .A1(n11999), .S(n3808), .Z(n12019) );
  CMXI2X1 U22281 ( .A0(n11988), .A1(n12019), .S(n3410), .Z(N5953) );
  CMX2X1 U22282 ( .A0(N7469), .A1(N7468), .S(n3869), .Z(n11995) );
  CMXI2X1 U22283 ( .A0(n11995), .A1(n11989), .S(n4086), .Z(n12009) );
  CMX2X1 U22284 ( .A0(n11990), .A1(n12009), .S(n3809), .Z(n12022) );
  CMXI2X1 U22285 ( .A0(n11991), .A1(n12022), .S(n3410), .Z(N5954) );
  CMX2X1 U22286 ( .A0(N7468), .A1(N7467), .S(n3863), .Z(n11998) );
  CMXI2X1 U22287 ( .A0(n11998), .A1(n11992), .S(n4086), .Z(n12012) );
  CMX2X1 U22288 ( .A0(n11993), .A1(n12012), .S(n3810), .Z(n12025) );
  CMXI2X1 U22289 ( .A0(n11994), .A1(n12025), .S(n3410), .Z(N5955) );
  CMX2X1 U22290 ( .A0(N7467), .A1(N7466), .S(n3864), .Z(n12008) );
  CMXI2X1 U22291 ( .A0(n12008), .A1(n11995), .S(n4086), .Z(n12015) );
  CMX2X1 U22292 ( .A0(n11996), .A1(n12015), .S(n3811), .Z(n12028) );
  CMXI2X1 U22293 ( .A0(n11997), .A1(n12028), .S(n3448), .Z(N5956) );
  CMX2X1 U22294 ( .A0(N7466), .A1(N7465), .S(n3880), .Z(n12011) );
  CMXI2X1 U22295 ( .A0(n12011), .A1(n11998), .S(n4086), .Z(n12018) );
  CMX2X1 U22296 ( .A0(n11999), .A1(n12018), .S(n3771), .Z(n12031) );
  CMXI2X1 U22297 ( .A0(n12000), .A1(n12031), .S(n3448), .Z(N5957) );
  CMXI2X1 U22298 ( .A0(n12071), .A1(n12001), .S(n4086), .Z(n12138) );
  CMX2X1 U22299 ( .A0(n12002), .A1(n12138), .S(n3807), .Z(n12273) );
  CMXI2X1 U22300 ( .A0(n12003), .A1(n12273), .S(n3448), .Z(N5237) );
  CMXI2X1 U22301 ( .A0(n4422), .A1(n12005), .S(n3799), .Z(n12007) );
  CMXI2X1 U22302 ( .A0(n12007), .A1(n12006), .S(n3448), .Z(N5165) );
  CMX2X1 U22303 ( .A0(N7465), .A1(N7464), .S(n3862), .Z(n12014) );
  CMXI2X1 U22304 ( .A0(n12014), .A1(n12008), .S(n4086), .Z(n12021) );
  CMX2X1 U22305 ( .A0(n12009), .A1(n12021), .S(n3808), .Z(n12034) );
  CMXI2X1 U22306 ( .A0(n12010), .A1(n12034), .S(n3447), .Z(N5958) );
  CMX2X1 U22307 ( .A0(N7464), .A1(N7463), .S(n3863), .Z(n12017) );
  CMXI2X1 U22308 ( .A0(n12017), .A1(n12011), .S(n4086), .Z(n12024) );
  CMX2X1 U22309 ( .A0(n12012), .A1(n12024), .S(n3809), .Z(n12037) );
  CMXI2X1 U22310 ( .A0(n12013), .A1(n12037), .S(n3447), .Z(N5959) );
  CMX2X1 U22311 ( .A0(N7463), .A1(N7462), .S(n3880), .Z(n12020) );
  CMXI2X1 U22312 ( .A0(n12020), .A1(n12014), .S(n4086), .Z(n12027) );
  CMX2X1 U22313 ( .A0(n12015), .A1(n12027), .S(n3810), .Z(n12043) );
  CMXI2X1 U22314 ( .A0(n12016), .A1(n12043), .S(n3447), .Z(N5960) );
  CMX2X1 U22315 ( .A0(N7462), .A1(N7461), .S(n3881), .Z(n12023) );
  CMXI2X1 U22316 ( .A0(n12023), .A1(n12017), .S(n4086), .Z(n12030) );
  CMX2X1 U22317 ( .A0(n12018), .A1(n12030), .S(n3811), .Z(n12046) );
  CMXI2X1 U22318 ( .A0(n12019), .A1(n12046), .S(n3447), .Z(N5961) );
  CMX2X1 U22319 ( .A0(N7461), .A1(N7460), .S(n3862), .Z(n12026) );
  CMXI2X1 U22320 ( .A0(n12026), .A1(n12020), .S(n4086), .Z(n12033) );
  CMX2X1 U22321 ( .A0(n12021), .A1(n12033), .S(n3812), .Z(n12049) );
  CMXI2X1 U22322 ( .A0(n12022), .A1(n12049), .S(n3447), .Z(N5962) );
  CMX2X1 U22323 ( .A0(N7460), .A1(N7459), .S(n3863), .Z(n12029) );
  CMXI2X1 U22324 ( .A0(n12029), .A1(n12023), .S(n4086), .Z(n12036) );
  CMX2X1 U22325 ( .A0(n12024), .A1(n12036), .S(n4316), .Z(n12052) );
  CMXI2X1 U22326 ( .A0(n12025), .A1(n12052), .S(n3447), .Z(N5963) );
  CMX2X1 U22327 ( .A0(N7459), .A1(N7458), .S(n3865), .Z(n12032) );
  CMXI2X1 U22328 ( .A0(n12032), .A1(n12026), .S(n4086), .Z(n12042) );
  CMX2X1 U22329 ( .A0(n12027), .A1(n12042), .S(n3771), .Z(n12055) );
  CMXI2X1 U22330 ( .A0(n12028), .A1(n12055), .S(n3447), .Z(N5964) );
  CMX2X1 U22331 ( .A0(N7458), .A1(N7457), .S(n3865), .Z(n12035) );
  CMXI2X1 U22332 ( .A0(n12035), .A1(n12029), .S(n4086), .Z(n12045) );
  CMX2X1 U22333 ( .A0(n12030), .A1(n12045), .S(n3772), .Z(n12058) );
  CMXI2X1 U22334 ( .A0(n12031), .A1(n12058), .S(n3447), .Z(N5965) );
  CMX2X1 U22335 ( .A0(N7457), .A1(N7456), .S(n3866), .Z(n12041) );
  CMXI2X1 U22336 ( .A0(n12041), .A1(n12032), .S(n4086), .Z(n12048) );
  CMX2X1 U22337 ( .A0(n12033), .A1(n12048), .S(n3773), .Z(n12061) );
  CMXI2X1 U22338 ( .A0(n12034), .A1(n12061), .S(n3447), .Z(N5966) );
  CMX2X1 U22339 ( .A0(N7456), .A1(N7455), .S(n3867), .Z(n12044) );
  CMXI2X1 U22340 ( .A0(n12044), .A1(n12035), .S(n4086), .Z(n12051) );
  CMX2X1 U22341 ( .A0(n12036), .A1(n12051), .S(n3774), .Z(n12064) );
  CMXI2X1 U22342 ( .A0(n12037), .A1(n12064), .S(n3447), .Z(N5967) );
  CMXI2X1 U22343 ( .A0(n12104), .A1(n12038), .S(n4085), .Z(n12171) );
  CMX2X1 U22344 ( .A0(n12039), .A1(n12171), .S(n3775), .Z(n12306) );
  CMXI2X1 U22345 ( .A0(n12040), .A1(n12306), .S(n3447), .Z(N5238) );
  CMX2X1 U22346 ( .A0(N7455), .A1(N7454), .S(n3869), .Z(n12047) );
  CMXI2X1 U22347 ( .A0(n12047), .A1(n12041), .S(n4085), .Z(n12054) );
  CMX2X1 U22348 ( .A0(n12042), .A1(n12054), .S(n3776), .Z(n12067) );
  CMXI2X1 U22349 ( .A0(n12043), .A1(n12067), .S(n3446), .Z(N5968) );
  CMX2X1 U22350 ( .A0(N7454), .A1(N7453), .S(n3870), .Z(n12050) );
  CMXI2X1 U22351 ( .A0(n12050), .A1(n12044), .S(n4085), .Z(n12057) );
  CMX2X1 U22352 ( .A0(n12045), .A1(n12057), .S(n3777), .Z(n12070) );
  CMXI2X1 U22353 ( .A0(n12046), .A1(n12070), .S(n3446), .Z(N5969) );
  CMX2X1 U22354 ( .A0(N7453), .A1(N7452), .S(n3871), .Z(n12053) );
  CMXI2X1 U22355 ( .A0(n12053), .A1(n12047), .S(n4085), .Z(n12060) );
  CMX2X1 U22356 ( .A0(n12048), .A1(n12060), .S(n3790), .Z(n12076) );
  CMXI2X1 U22357 ( .A0(n12049), .A1(n12076), .S(n3446), .Z(N5970) );
  CMX2X1 U22358 ( .A0(N7452), .A1(N7451), .S(n3870), .Z(n12056) );
  CMXI2X1 U22359 ( .A0(n12056), .A1(n12050), .S(n4085), .Z(n12063) );
  CMX2X1 U22360 ( .A0(n12051), .A1(n12063), .S(n3791), .Z(n12079) );
  CMXI2X1 U22361 ( .A0(n12052), .A1(n12079), .S(n3449), .Z(N5971) );
  CMX2X1 U22362 ( .A0(N7451), .A1(N7450), .S(n3871), .Z(n12059) );
  CMXI2X1 U22363 ( .A0(n12059), .A1(n12053), .S(n4085), .Z(n12066) );
  CMX2X1 U22364 ( .A0(n12054), .A1(n12066), .S(n3794), .Z(n12082) );
  CMXI2X1 U22365 ( .A0(n12055), .A1(n12082), .S(n3449), .Z(N5972) );
  CMX2X1 U22366 ( .A0(N7450), .A1(N7449), .S(n3872), .Z(n12062) );
  CMXI2X1 U22367 ( .A0(n12062), .A1(n12056), .S(n4085), .Z(n12069) );
  CMX2X1 U22368 ( .A0(n12057), .A1(n12069), .S(n3795), .Z(n12085) );
  CMXI2X1 U22369 ( .A0(n12058), .A1(n12085), .S(n3449), .Z(N5973) );
  CMX2X1 U22370 ( .A0(N7449), .A1(N7448), .S(n3873), .Z(n12065) );
  CMXI2X1 U22371 ( .A0(n12065), .A1(n12059), .S(n4085), .Z(n12075) );
  CMX2X1 U22372 ( .A0(n12060), .A1(n12075), .S(n3812), .Z(n12088) );
  CMXI2X1 U22373 ( .A0(n12061), .A1(n12088), .S(n3449), .Z(N5974) );
  CMX2X1 U22374 ( .A0(N7448), .A1(N7447), .S(n3864), .Z(n12068) );
  CMXI2X1 U22375 ( .A0(n12068), .A1(n12062), .S(n4085), .Z(n12078) );
  CMX2X1 U22376 ( .A0(n12063), .A1(n12078), .S(n4313), .Z(n12091) );
  CMXI2X1 U22377 ( .A0(n12064), .A1(n12091), .S(n3449), .Z(N5975) );
  CMX2X1 U22378 ( .A0(N7447), .A1(N7446), .S(n3865), .Z(n12074) );
  CMXI2X1 U22379 ( .A0(n12074), .A1(n12065), .S(n4085), .Z(n12081) );
  CMX2X1 U22380 ( .A0(n12066), .A1(n12081), .S(n3771), .Z(n12094) );
  CMXI2X1 U22381 ( .A0(n12067), .A1(n12094), .S(n3449), .Z(N5976) );
  CMX2X1 U22382 ( .A0(N7446), .A1(N7445), .S(n3866), .Z(n12077) );
  CMXI2X1 U22383 ( .A0(n12077), .A1(n12068), .S(n4085), .Z(n12084) );
  CMX2X1 U22384 ( .A0(n12069), .A1(n12084), .S(n3772), .Z(n12097) );
  CMXI2X1 U22385 ( .A0(n12070), .A1(n12097), .S(n3449), .Z(N5977) );
  CMX2X1 U22386 ( .A0(N8184), .A1(N8183), .S(n3867), .Z(n12137) );
  CMXI2X1 U22387 ( .A0(n12137), .A1(n12071), .S(n4085), .Z(n12204) );
  CMX2X1 U22388 ( .A0(n12072), .A1(n12204), .S(n3773), .Z(n12339) );
  CMXI2X1 U22389 ( .A0(n12073), .A1(n12339), .S(n3449), .Z(N5239) );
  CMX2X1 U22390 ( .A0(N7445), .A1(N7444), .S(n3864), .Z(n12080) );
  CMXI2X1 U22391 ( .A0(n12080), .A1(n12074), .S(n4085), .Z(n12087) );
  CMX2X1 U22392 ( .A0(n12075), .A1(n12087), .S(n3772), .Z(n12100) );
  CMXI2X1 U22393 ( .A0(n12076), .A1(n12100), .S(n3449), .Z(N5978) );
  CMX2X1 U22394 ( .A0(N7444), .A1(N7443), .S(n3877), .Z(n12083) );
  CMXI2X1 U22395 ( .A0(n12083), .A1(n12077), .S(n4085), .Z(n12090) );
  CMX2X1 U22396 ( .A0(n12078), .A1(n12090), .S(n3792), .Z(n12103) );
  CMXI2X1 U22397 ( .A0(n12079), .A1(n12103), .S(n3449), .Z(N5979) );
  CMX2X1 U22398 ( .A0(N7443), .A1(N7442), .S(n3878), .Z(n12086) );
  CMXI2X1 U22399 ( .A0(n12086), .A1(n12080), .S(n4085), .Z(n12093) );
  CMX2X1 U22400 ( .A0(n12081), .A1(n12093), .S(n3793), .Z(n12109) );
  CMXI2X1 U22401 ( .A0(n12082), .A1(n12109), .S(n3449), .Z(N5980) );
  CMX2X1 U22402 ( .A0(N7442), .A1(N7441), .S(n3862), .Z(n12089) );
  CMXI2X1 U22403 ( .A0(n12089), .A1(n12083), .S(n4085), .Z(n12096) );
  CMX2X1 U22404 ( .A0(n12084), .A1(n12096), .S(n3794), .Z(n12112) );
  CMXI2X1 U22405 ( .A0(n12085), .A1(n12112), .S(n3448), .Z(N5981) );
  CMX2X1 U22406 ( .A0(N7441), .A1(N7440), .S(n3863), .Z(n12092) );
  CMXI2X1 U22407 ( .A0(n12092), .A1(n12086), .S(n4084), .Z(n12099) );
  CMX2X1 U22408 ( .A0(n12087), .A1(n12099), .S(n3795), .Z(n12115) );
  CMXI2X1 U22409 ( .A0(n12088), .A1(n12115), .S(n3448), .Z(N5982) );
  CMX2X1 U22410 ( .A0(N7440), .A1(N7439), .S(n3864), .Z(n12095) );
  CMXI2X1 U22411 ( .A0(n12095), .A1(n12089), .S(n4084), .Z(n12102) );
  CMX2X1 U22412 ( .A0(n12090), .A1(n12102), .S(n3796), .Z(n12118) );
  CMXI2X1 U22413 ( .A0(n12091), .A1(n12118), .S(n3448), .Z(N5983) );
  CMX2X1 U22414 ( .A0(N7439), .A1(N7438), .S(n3865), .Z(n12098) );
  CMXI2X1 U22415 ( .A0(n12098), .A1(n12092), .S(n4084), .Z(n12108) );
  CMX2X1 U22416 ( .A0(n12093), .A1(n12108), .S(n3797), .Z(n12121) );
  CMXI2X1 U22417 ( .A0(n12094), .A1(n12121), .S(n3448), .Z(N5984) );
  CMX2X1 U22418 ( .A0(N7438), .A1(N7437), .S(n3866), .Z(n12101) );
  CMXI2X1 U22419 ( .A0(n12101), .A1(n12095), .S(n4084), .Z(n12111) );
  CMX2X1 U22420 ( .A0(n12096), .A1(n12111), .S(n3805), .Z(n12124) );
  CMXI2X1 U22421 ( .A0(n12097), .A1(n12124), .S(n3448), .Z(N5985) );
  CMX2X1 U22422 ( .A0(N7437), .A1(N7436), .S(n3867), .Z(n12107) );
  CMXI2X1 U22423 ( .A0(n12107), .A1(n12098), .S(n4084), .Z(n12114) );
  CMX2X1 U22424 ( .A0(n12099), .A1(n12114), .S(n3806), .Z(n12127) );
  CMXI2X1 U22425 ( .A0(n12100), .A1(n12127), .S(n3448), .Z(N5986) );
  CMX2X1 U22426 ( .A0(N7436), .A1(N7435), .S(n3868), .Z(n12110) );
  CMXI2X1 U22427 ( .A0(n12110), .A1(n12101), .S(n4084), .Z(n12117) );
  CMX2X1 U22428 ( .A0(n12102), .A1(n12117), .S(n3807), .Z(n12130) );
  CMXI2X1 U22429 ( .A0(n12103), .A1(n12130), .S(n3448), .Z(N5987) );
  CMXI2X1 U22430 ( .A0(n12170), .A1(n12104), .S(n4084), .Z(n12238) );
  CMX2X1 U22431 ( .A0(n12105), .A1(n12238), .S(n3808), .Z(n12374) );
  CMXI2X1 U22432 ( .A0(n12106), .A1(n12374), .S(n3451), .Z(N5240) );
  CMX2X1 U22433 ( .A0(N7435), .A1(N7434), .S(n3879), .Z(n12113) );
  CMXI2X1 U22434 ( .A0(n12113), .A1(n12107), .S(n4084), .Z(n12120) );
  CMX2X1 U22435 ( .A0(n12108), .A1(n12120), .S(n3809), .Z(n12133) );
  CMXI2X1 U22436 ( .A0(n12109), .A1(n12133), .S(n3451), .Z(N5988) );
  CMX2X1 U22437 ( .A0(N7434), .A1(N7433), .S(n3879), .Z(n12116) );
  CMXI2X1 U22438 ( .A0(n12116), .A1(n12110), .S(n4084), .Z(n12123) );
  CMX2X1 U22439 ( .A0(n12111), .A1(n12123), .S(n3810), .Z(n12136) );
  CMXI2X1 U22440 ( .A0(n12112), .A1(n12136), .S(n3451), .Z(N5989) );
  CMX2X1 U22441 ( .A0(N7433), .A1(N7432), .S(n3880), .Z(n12119) );
  CMXI2X1 U22442 ( .A0(n12119), .A1(n12113), .S(n4084), .Z(n12126) );
  CMX2X1 U22443 ( .A0(n12114), .A1(n12126), .S(n3811), .Z(n12142) );
  CMXI2X1 U22444 ( .A0(n12115), .A1(n12142), .S(n3451), .Z(N5990) );
  CMX2X1 U22445 ( .A0(N7432), .A1(N7431), .S(n3881), .Z(n12122) );
  CMXI2X1 U22446 ( .A0(n12122), .A1(n12116), .S(n4084), .Z(n12129) );
  CMX2X1 U22447 ( .A0(n12117), .A1(n12129), .S(n3812), .Z(n12145) );
  CMXI2X1 U22448 ( .A0(n12118), .A1(n12145), .S(n3451), .Z(N5991) );
  CMX2X1 U22449 ( .A0(N7431), .A1(N7430), .S(n3862), .Z(n12125) );
  CMXI2X1 U22450 ( .A0(n12125), .A1(n12119), .S(n4084), .Z(n12132) );
  CMX2X1 U22451 ( .A0(n12120), .A1(n12132), .S(n4315), .Z(n12148) );
  CMXI2X1 U22452 ( .A0(n12121), .A1(n12148), .S(n3451), .Z(N5992) );
  CMX2X1 U22453 ( .A0(N7430), .A1(N7429), .S(n3863), .Z(n12128) );
  CMXI2X1 U22454 ( .A0(n12128), .A1(n12122), .S(n4084), .Z(n12135) );
  CMX2X1 U22455 ( .A0(n12123), .A1(n12135), .S(n3771), .Z(n12151) );
  CMXI2X1 U22456 ( .A0(n12124), .A1(n12151), .S(n3451), .Z(N5993) );
  CMX2X1 U22457 ( .A0(N7429), .A1(N7428), .S(n3864), .Z(n12131) );
  CMXI2X1 U22458 ( .A0(n12131), .A1(n12125), .S(n4084), .Z(n12141) );
  CMX2X1 U22459 ( .A0(n12126), .A1(n12141), .S(n3795), .Z(n12154) );
  CMXI2X1 U22460 ( .A0(n12127), .A1(n12154), .S(n3450), .Z(N5994) );
  CMX2X1 U22461 ( .A0(N7428), .A1(N7427), .S(n3865), .Z(n12134) );
  CMXI2X1 U22462 ( .A0(n12134), .A1(n12128), .S(n4084), .Z(n12144) );
  CMX2X1 U22463 ( .A0(n12129), .A1(n12144), .S(n3796), .Z(n12157) );
  CMXI2X1 U22464 ( .A0(n12130), .A1(n12157), .S(n3450), .Z(N5995) );
  CMX2X1 U22465 ( .A0(N7427), .A1(N7426), .S(n3862), .Z(n12140) );
  CMXI2X1 U22466 ( .A0(n12140), .A1(n12131), .S(n4084), .Z(n12147) );
  CMX2X1 U22467 ( .A0(n12132), .A1(n12147), .S(n3774), .Z(n12160) );
  CMXI2X1 U22468 ( .A0(n12133), .A1(n12160), .S(n3450), .Z(N5996) );
  CMX2X1 U22469 ( .A0(N7426), .A1(N7425), .S(n3863), .Z(n12143) );
  CMXI2X1 U22470 ( .A0(n12143), .A1(n12134), .S(n4083), .Z(n12150) );
  CMX2X1 U22471 ( .A0(n12135), .A1(n12150), .S(n3775), .Z(n12163) );
  CMXI2X1 U22472 ( .A0(n12136), .A1(n12163), .S(n3450), .Z(N5997) );
  CMXI2X1 U22473 ( .A0(n12203), .A1(n12137), .S(n4083), .Z(n12272) );
  CMX2X1 U22474 ( .A0(n12138), .A1(n12272), .S(n3776), .Z(n12407) );
  CMXI2X1 U22475 ( .A0(n12139), .A1(n12407), .S(n3450), .Z(N5241) );
  CMX2X1 U22476 ( .A0(N7425), .A1(N7424), .S(n3867), .Z(n12146) );
  CMXI2X1 U22477 ( .A0(n12146), .A1(n12140), .S(n4083), .Z(n12153) );
  CMX2X1 U22478 ( .A0(n12141), .A1(n12153), .S(n3777), .Z(n12166) );
  CMXI2X1 U22479 ( .A0(n12142), .A1(n12166), .S(n3450), .Z(N5998) );
  CMX2X1 U22480 ( .A0(N7424), .A1(N7423), .S(n3865), .Z(n12149) );
  CMXI2X1 U22481 ( .A0(n12149), .A1(n12143), .S(n4083), .Z(n12156) );
  CMX2X1 U22482 ( .A0(n12144), .A1(n12156), .S(n3790), .Z(n12169) );
  CMX2X1 U22483 ( .A0(N7423), .A1(N7422), .S(n3866), .Z(n12152) );
  CMXI2X1 U22484 ( .A0(n12152), .A1(n12146), .S(n4083), .Z(n12159) );
  CMX2X1 U22485 ( .A0(n12147), .A1(n12159), .S(n3773), .Z(n12175) );
  CMXI2X1 U22486 ( .A0(n12148), .A1(n12175), .S(n3450), .Z(N6000) );
  CMX2X1 U22487 ( .A0(N7422), .A1(N7421), .S(n3867), .Z(n12155) );
  CMXI2X1 U22488 ( .A0(n12155), .A1(n12149), .S(n4083), .Z(n12162) );
  CMX2X1 U22489 ( .A0(n12150), .A1(n12162), .S(n3772), .Z(n12178) );
  CMXI2X1 U22490 ( .A0(n12151), .A1(n12178), .S(n3450), .Z(N6001) );
  CMX2X1 U22491 ( .A0(N7421), .A1(N7420), .S(n3866), .Z(n12158) );
  CMXI2X1 U22492 ( .A0(n12158), .A1(n12152), .S(n4083), .Z(n12165) );
  CMX2X1 U22493 ( .A0(n12153), .A1(n12165), .S(n3773), .Z(n12181) );
  CMXI2X1 U22494 ( .A0(n12154), .A1(n12181), .S(n3450), .Z(N6002) );
  CMX2X1 U22495 ( .A0(N7420), .A1(N7419), .S(n3874), .Z(n12161) );
  CMXI2X1 U22496 ( .A0(n12161), .A1(n12155), .S(n4083), .Z(n12168) );
  CMX2X1 U22497 ( .A0(n12156), .A1(n12168), .S(n3774), .Z(n12184) );
  CMXI2X1 U22498 ( .A0(n12157), .A1(n12184), .S(n3450), .Z(N6003) );
  CMX2X1 U22499 ( .A0(N7419), .A1(N7418), .S(n3875), .Z(n12164) );
  CMXI2X1 U22500 ( .A0(n12164), .A1(n12158), .S(n4083), .Z(n12174) );
  CMX2X1 U22501 ( .A0(n12159), .A1(n12174), .S(n3775), .Z(n12187) );
  CMXI2X1 U22502 ( .A0(n12160), .A1(n12187), .S(n3453), .Z(N6004) );
  CMX2X1 U22503 ( .A0(N7418), .A1(N7417), .S(n3876), .Z(n12167) );
  CMXI2X1 U22504 ( .A0(n12167), .A1(n12161), .S(n4083), .Z(n12177) );
  CMX2X1 U22505 ( .A0(n12162), .A1(n12177), .S(n3776), .Z(n12190) );
  CMXI2X1 U22506 ( .A0(n12163), .A1(n12190), .S(n3453), .Z(N6005) );
  CMX2X1 U22507 ( .A0(N7417), .A1(N7416), .S(n3877), .Z(n12173) );
  CMXI2X1 U22508 ( .A0(n12173), .A1(n12164), .S(n4083), .Z(n12180) );
  CMX2X1 U22509 ( .A0(n12165), .A1(n12180), .S(n3777), .Z(n12193) );
  CMXI2X1 U22510 ( .A0(n12166), .A1(n12193), .S(n3453), .Z(N6006) );
  CMX2X1 U22511 ( .A0(N7416), .A1(N7415), .S(n3878), .Z(n12176) );
  CMXI2X1 U22512 ( .A0(n12176), .A1(n12167), .S(n4083), .Z(n12183) );
  CMX2X1 U22513 ( .A0(n12168), .A1(n12183), .S(n3790), .Z(n12196) );
  CMXI2X1 U22514 ( .A0(n12236), .A1(n12170), .S(n4083), .Z(n12305) );
  CMX2X1 U22515 ( .A0(n12171), .A1(n12305), .S(n3791), .Z(n12439) );
  CMXI2X1 U22516 ( .A0(n12172), .A1(n12439), .S(n3452), .Z(N5242) );
  CMX2X1 U22517 ( .A0(N7415), .A1(N7414), .S(n3880), .Z(n12179) );
  CMXI2X1 U22518 ( .A0(n12179), .A1(n12173), .S(n4083), .Z(n12186) );
  CMX2X1 U22519 ( .A0(n12174), .A1(n12186), .S(n3792), .Z(n12199) );
  CMXI2X1 U22520 ( .A0(n12175), .A1(n12199), .S(n3452), .Z(N6008) );
  CMX2X1 U22521 ( .A0(N7414), .A1(N7413), .S(n3872), .Z(n12182) );
  CMXI2X1 U22522 ( .A0(n12182), .A1(n12176), .S(n4083), .Z(n12189) );
  CMX2X1 U22523 ( .A0(n12177), .A1(n12189), .S(n3793), .Z(n12202) );
  CMXI2X1 U22524 ( .A0(n12178), .A1(n12202), .S(n3452), .Z(N6009) );
  CMX2X1 U22525 ( .A0(N7413), .A1(N7412), .S(n3873), .Z(n12185) );
  CMXI2X1 U22526 ( .A0(n12185), .A1(n12179), .S(n4083), .Z(n12192) );
  CMX2X1 U22527 ( .A0(n12180), .A1(n12192), .S(n3794), .Z(n12208) );
  CMXI2X1 U22528 ( .A0(n12181), .A1(n12208), .S(n3452), .Z(N6010) );
  CMX2X1 U22529 ( .A0(N7412), .A1(N7411), .S(n3881), .Z(n12188) );
  CMXI2X1 U22530 ( .A0(n12188), .A1(n12182), .S(n4082), .Z(n12195) );
  CMX2X1 U22531 ( .A0(n12183), .A1(n12195), .S(n3795), .Z(n12211) );
  CMXI2X1 U22532 ( .A0(n12184), .A1(n12211), .S(n3452), .Z(N6011) );
  CMX2X1 U22533 ( .A0(N7411), .A1(N7410), .S(n3862), .Z(n12191) );
  CMXI2X1 U22534 ( .A0(n12191), .A1(n12185), .S(n4082), .Z(n12198) );
  CMX2X1 U22535 ( .A0(n12186), .A1(n12198), .S(n3796), .Z(n12214) );
  CMXI2X1 U22536 ( .A0(n12187), .A1(n12214), .S(n3452), .Z(N6012) );
  CMX2X1 U22537 ( .A0(N7410), .A1(N7409), .S(n3868), .Z(n12194) );
  CMXI2X1 U22538 ( .A0(n12194), .A1(n12188), .S(n4082), .Z(n12201) );
  CMX2X1 U22539 ( .A0(n12189), .A1(n12201), .S(n3797), .Z(n12217) );
  CMXI2X1 U22540 ( .A0(n12190), .A1(n12217), .S(n3452), .Z(N6013) );
  CMX2X1 U22541 ( .A0(N7409), .A1(N7408), .S(n3869), .Z(n12197) );
  CMXI2X1 U22542 ( .A0(n12197), .A1(n12191), .S(n4082), .Z(n12207) );
  CMX2X1 U22543 ( .A0(n12192), .A1(n12207), .S(n3805), .Z(n12220) );
  CMXI2X1 U22544 ( .A0(n12193), .A1(n12220), .S(n3452), .Z(N6014) );
  CMX2X1 U22545 ( .A0(N7408), .A1(N7407), .S(n3870), .Z(n12200) );
  CMXI2X1 U22546 ( .A0(n12200), .A1(n12194), .S(n4082), .Z(n12210) );
  CMX2X1 U22547 ( .A0(n12195), .A1(n12210), .S(n3806), .Z(n12223) );
  CMXI2X1 U22548 ( .A0(n12196), .A1(n12223), .S(n3452), .Z(N6015) );
  CMX2X1 U22549 ( .A0(N7407), .A1(N7406), .S(n3871), .Z(n12206) );
  CMXI2X1 U22550 ( .A0(n12206), .A1(n12197), .S(n4082), .Z(n12213) );
  CMX2X1 U22551 ( .A0(n12198), .A1(n12213), .S(n3796), .Z(n12226) );
  CMXI2X1 U22552 ( .A0(n12199), .A1(n12226), .S(n3452), .Z(N6016) );
  CMX2X1 U22553 ( .A0(N7406), .A1(N7405), .S(n3869), .Z(n12209) );
  CMXI2X1 U22554 ( .A0(n12209), .A1(n12200), .S(n4082), .Z(n12216) );
  CMX2X1 U22555 ( .A0(n12201), .A1(n12216), .S(n3795), .Z(n12229) );
  CMXI2X1 U22556 ( .A0(n12202), .A1(n12229), .S(n3451), .Z(N6017) );
  CMXI2X1 U22557 ( .A0(n12270), .A1(n12203), .S(n4082), .Z(n12338) );
  CMX2X1 U22558 ( .A0(n12204), .A1(n12338), .S(n3796), .Z(n12471) );
  CMXI2X1 U22559 ( .A0(n12205), .A1(n12471), .S(n3451), .Z(N5243) );
  CMX2X1 U22560 ( .A0(N7405), .A1(N7404), .S(n3879), .Z(n12212) );
  CMXI2X1 U22561 ( .A0(n12212), .A1(n12206), .S(n4082), .Z(n12219) );
  CMX2X1 U22562 ( .A0(n12207), .A1(n12219), .S(n3797), .Z(n12232) );
  CMXI2X1 U22563 ( .A0(n12208), .A1(n12232), .S(n3451), .Z(N6018) );
  CMX2X1 U22564 ( .A0(N7404), .A1(N7403), .S(n3880), .Z(n12215) );
  CMXI2X1 U22565 ( .A0(n12215), .A1(n12209), .S(n4082), .Z(n12222) );
  CMX2X1 U22566 ( .A0(n12210), .A1(n12222), .S(n3805), .Z(n12235) );
  CMXI2X1 U22567 ( .A0(n12211), .A1(n12235), .S(n3451), .Z(N6019) );
  CMX2X1 U22568 ( .A0(N7403), .A1(N7402), .S(n3881), .Z(n12218) );
  CMXI2X1 U22569 ( .A0(n12218), .A1(n12212), .S(n4082), .Z(n12225) );
  CMX2X1 U22570 ( .A0(n12213), .A1(n12225), .S(n3806), .Z(n12242) );
  CMXI2X1 U22571 ( .A0(n12214), .A1(n12242), .S(n3454), .Z(N6020) );
  CMX2X1 U22572 ( .A0(N7402), .A1(N7401), .S(n3870), .Z(n12221) );
  CMXI2X1 U22573 ( .A0(n12221), .A1(n12215), .S(n4082), .Z(n12228) );
  CMX2X1 U22574 ( .A0(n12216), .A1(n12228), .S(n3807), .Z(n12245) );
  CMXI2X1 U22575 ( .A0(n12217), .A1(n12245), .S(n3454), .Z(N6021) );
  CMX2X1 U22576 ( .A0(N7401), .A1(N7400), .S(n3871), .Z(n12224) );
  CMXI2X1 U22577 ( .A0(n12224), .A1(n12218), .S(n4082), .Z(n12231) );
  CMX2X1 U22578 ( .A0(n12219), .A1(n12231), .S(n3808), .Z(n12248) );
  CMXI2X1 U22579 ( .A0(n12220), .A1(n12248), .S(n3454), .Z(N6022) );
  CMX2X1 U22580 ( .A0(N7400), .A1(N7399), .S(n3862), .Z(n12227) );
  CMXI2X1 U22581 ( .A0(n12227), .A1(n12221), .S(n4082), .Z(n12234) );
  CMX2X1 U22582 ( .A0(n12222), .A1(n12234), .S(n3809), .Z(n12251) );
  CMXI2X1 U22583 ( .A0(n12223), .A1(n12251), .S(n3454), .Z(N6023) );
  CMX2X1 U22584 ( .A0(N7399), .A1(N7398), .S(n3863), .Z(n12230) );
  CMXI2X1 U22585 ( .A0(n12230), .A1(n12224), .S(n4082), .Z(n12241) );
  CMX2X1 U22586 ( .A0(n12225), .A1(n12241), .S(n3810), .Z(n12254) );
  CMXI2X1 U22587 ( .A0(n12226), .A1(n12254), .S(n3454), .Z(N6024) );
  CMX2X1 U22588 ( .A0(N7398), .A1(N7397), .S(n3872), .Z(n12233) );
  CMXI2X1 U22589 ( .A0(n12233), .A1(n12227), .S(n4082), .Z(n12244) );
  CMX2X1 U22590 ( .A0(n12228), .A1(n12244), .S(n3811), .Z(n12257) );
  CMXI2X1 U22591 ( .A0(n12229), .A1(n12257), .S(n3454), .Z(N6025) );
  CMX2X1 U22592 ( .A0(N7397), .A1(N7396), .S(n3873), .Z(n12240) );
  CMXI2X1 U22593 ( .A0(n12240), .A1(n12230), .S(n4081), .Z(n12247) );
  CMX2X1 U22594 ( .A0(n12231), .A1(n12247), .S(n3812), .Z(n12260) );
  CMXI2X1 U22595 ( .A0(n12232), .A1(n12260), .S(n3454), .Z(N6026) );
  CMX2X1 U22596 ( .A0(N7396), .A1(N7395), .S(n3874), .Z(n12243) );
  CMXI2X1 U22597 ( .A0(n12243), .A1(n12233), .S(n4081), .Z(n12250) );
  CMX2X1 U22598 ( .A0(n12234), .A1(n12250), .S(n4309), .Z(n12263) );
  CMXI2X1 U22599 ( .A0(n12235), .A1(n12263), .S(n3454), .Z(N6027) );
  CMXI2X1 U22600 ( .A0(n12237), .A1(n12236), .S(n4081), .Z(n12373) );
  CMX2X1 U22601 ( .A0(n12238), .A1(n12373), .S(n3790), .Z(n12503) );
  CMXI2X1 U22602 ( .A0(n12239), .A1(n12503), .S(n3454), .Z(N5244) );
  CMX2X1 U22603 ( .A0(N7395), .A1(N7394), .S(n3875), .Z(n12246) );
  CMXI2X1 U22604 ( .A0(n12246), .A1(n12240), .S(n4081), .Z(n12253) );
  CMX2X1 U22605 ( .A0(n12241), .A1(n12253), .S(n3772), .Z(n12266) );
  CMXI2X1 U22606 ( .A0(n12242), .A1(n12266), .S(n3454), .Z(N6028) );
  CMX2X1 U22607 ( .A0(N7394), .A1(N7393), .S(n3876), .Z(n12249) );
  CMXI2X1 U22608 ( .A0(n12249), .A1(n12243), .S(n4081), .Z(n12256) );
  CMX2X1 U22609 ( .A0(n12244), .A1(n12256), .S(n3773), .Z(n12269) );
  CMXI2X1 U22610 ( .A0(n12245), .A1(n12269), .S(n3453), .Z(N6029) );
  CMX2X1 U22611 ( .A0(N7393), .A1(N7392), .S(n3877), .Z(n12252) );
  CMXI2X1 U22612 ( .A0(n12252), .A1(n12246), .S(n4081), .Z(n12259) );
  CMX2X1 U22613 ( .A0(n12247), .A1(n12259), .S(n3774), .Z(n12276) );
  CMXI2X1 U22614 ( .A0(n12248), .A1(n12276), .S(n3453), .Z(N6030) );
  CMX2X1 U22615 ( .A0(N7392), .A1(N7391), .S(n3881), .Z(n12255) );
  CMXI2X1 U22616 ( .A0(n12255), .A1(n12249), .S(n4081), .Z(n12262) );
  CMX2X1 U22617 ( .A0(n12250), .A1(n12262), .S(n3775), .Z(n12279) );
  CMXI2X1 U22618 ( .A0(n12251), .A1(n12279), .S(n3453), .Z(N6031) );
  CMX2X1 U22619 ( .A0(N7391), .A1(N7390), .S(n3877), .Z(n12258) );
  CMXI2X1 U22620 ( .A0(n12258), .A1(n12252), .S(n4081), .Z(n12265) );
  CMX2X1 U22621 ( .A0(n12253), .A1(n12265), .S(n3776), .Z(n12282) );
  CMXI2X1 U22622 ( .A0(n12254), .A1(n12282), .S(n3453), .Z(N6032) );
  CMX2X1 U22623 ( .A0(N7390), .A1(N7389), .S(n3878), .Z(n12261) );
  CMXI2X1 U22624 ( .A0(n12261), .A1(n12255), .S(n4081), .Z(n12268) );
  CMX2X1 U22625 ( .A0(n12256), .A1(n12268), .S(n3777), .Z(n12285) );
  CMXI2X1 U22626 ( .A0(n12257), .A1(n12285), .S(n3453), .Z(N6033) );
  CMX2X1 U22627 ( .A0(N7389), .A1(N7388), .S(n3879), .Z(n12264) );
  CMXI2X1 U22628 ( .A0(n12264), .A1(n12258), .S(n4081), .Z(n12275) );
  CMX2X1 U22629 ( .A0(n12259), .A1(n12275), .S(n3790), .Z(n12288) );
  CMXI2X1 U22630 ( .A0(n12260), .A1(n12288), .S(n3453), .Z(N6034) );
  CMX2X1 U22631 ( .A0(N7388), .A1(N7387), .S(n3880), .Z(n12267) );
  CMXI2X1 U22632 ( .A0(n12267), .A1(n12261), .S(n4081), .Z(n12278) );
  CMX2X1 U22633 ( .A0(n12262), .A1(n12278), .S(n3791), .Z(n12291) );
  CMXI2X1 U22634 ( .A0(n12263), .A1(n12291), .S(n3453), .Z(N6035) );
  CMX2X1 U22635 ( .A0(N7387), .A1(N7386), .S(n3881), .Z(n12274) );
  CMXI2X1 U22636 ( .A0(n12274), .A1(n12264), .S(n4081), .Z(n12281) );
  CMX2X1 U22637 ( .A0(n12265), .A1(n12281), .S(n3792), .Z(n12294) );
  CMXI2X1 U22638 ( .A0(n12266), .A1(n12294), .S(n3453), .Z(N6036) );
  CMX2X1 U22639 ( .A0(N7386), .A1(N7385), .S(n3862), .Z(n12277) );
  CMXI2X1 U22640 ( .A0(n12277), .A1(n12267), .S(n4081), .Z(n12284) );
  CMX2X1 U22641 ( .A0(n12268), .A1(n12284), .S(n3793), .Z(n12297) );
  CMXI2X1 U22642 ( .A0(n12269), .A1(n12297), .S(n3443), .Z(N6037) );
  CMXI2X1 U22643 ( .A0(n12271), .A1(n12270), .S(n4081), .Z(n12406) );
  CMX2X1 U22644 ( .A0(n12272), .A1(n12406), .S(n3794), .Z(n12535) );
  CMXI2X1 U22645 ( .A0(n12273), .A1(n12535), .S(n3274), .Z(N5245) );
  CMX2X1 U22646 ( .A0(N7385), .A1(N7384), .S(n3863), .Z(n12280) );
  CMXI2X1 U22647 ( .A0(n12280), .A1(n12274), .S(n4081), .Z(n12287) );
  CMX2X1 U22648 ( .A0(n12275), .A1(n12287), .S(n3795), .Z(n12300) );
  CMXI2X1 U22649 ( .A0(n12276), .A1(n12300), .S(n3274), .Z(N6038) );
  CMX2X1 U22650 ( .A0(N7384), .A1(N7383), .S(n3866), .Z(n12283) );
  CMXI2X1 U22651 ( .A0(n12283), .A1(n12277), .S(n4081), .Z(n12290) );
  CMX2X1 U22652 ( .A0(n12278), .A1(n12290), .S(n3796), .Z(n12303) );
  CMXI2X1 U22653 ( .A0(n12279), .A1(n12303), .S(n3274), .Z(N6039) );
  CMX2X1 U22654 ( .A0(N7383), .A1(N7382), .S(n3867), .Z(n12286) );
  CMXI2X1 U22655 ( .A0(n12286), .A1(n12280), .S(n4080), .Z(n12293) );
  CMX2X1 U22656 ( .A0(n12281), .A1(n12293), .S(n3797), .Z(n12309) );
  CMXI2X1 U22657 ( .A0(n12282), .A1(n12309), .S(n3274), .Z(N6040) );
  CMX2X1 U22658 ( .A0(N7382), .A1(N7381), .S(n3864), .Z(n12289) );
  CMXI2X1 U22659 ( .A0(n12289), .A1(n12283), .S(n4080), .Z(n12296) );
  CMX2X1 U22660 ( .A0(n12284), .A1(n12296), .S(n3805), .Z(n12312) );
  CMXI2X1 U22661 ( .A0(n12285), .A1(n12312), .S(n3274), .Z(N6041) );
  CMX2X1 U22662 ( .A0(N7381), .A1(N7380), .S(n3865), .Z(n12292) );
  CMXI2X1 U22663 ( .A0(n12292), .A1(n12286), .S(n4080), .Z(n12299) );
  CMX2X1 U22664 ( .A0(n12287), .A1(n12299), .S(n3806), .Z(n12315) );
  CMXI2X1 U22665 ( .A0(n12288), .A1(n12315), .S(n3274), .Z(N6042) );
  CMX2X1 U22666 ( .A0(N7380), .A1(N7379), .S(n3874), .Z(n12295) );
  CMXI2X1 U22667 ( .A0(n12295), .A1(n12289), .S(n4080), .Z(n12302) );
  CMX2X1 U22668 ( .A0(n12290), .A1(n12302), .S(n3772), .Z(n12318) );
  CMXI2X1 U22669 ( .A0(n12291), .A1(n12318), .S(n3274), .Z(N6043) );
  CMX2X1 U22670 ( .A0(N7379), .A1(N7378), .S(n3875), .Z(n12298) );
  CMXI2X1 U22671 ( .A0(n12298), .A1(n12292), .S(n4080), .Z(n12308) );
  CMX2X1 U22672 ( .A0(n12293), .A1(n12308), .S(n3773), .Z(n12321) );
  CMXI2X1 U22673 ( .A0(n12294), .A1(n12321), .S(n3274), .Z(N6044) );
  CMX2X1 U22674 ( .A0(N7378), .A1(N7377), .S(n3876), .Z(n12301) );
  CMXI2X1 U22675 ( .A0(n12301), .A1(n12295), .S(n4080), .Z(n12311) );
  CMX2X1 U22676 ( .A0(n12296), .A1(n12311), .S(n3810), .Z(n12324) );
  CMXI2X1 U22677 ( .A0(n12297), .A1(n12324), .S(n3274), .Z(N6045) );
  CMX2X1 U22678 ( .A0(N7377), .A1(N7376), .S(n3877), .Z(n12307) );
  CMXI2X1 U22679 ( .A0(n12307), .A1(n12298), .S(n4080), .Z(n12314) );
  CMX2X1 U22680 ( .A0(n12299), .A1(n12314), .S(n3811), .Z(n12327) );
  CMXI2X1 U22681 ( .A0(n12300), .A1(n12327), .S(n3274), .Z(N6046) );
  CMX2X1 U22682 ( .A0(N7376), .A1(N7375), .S(n3864), .Z(n12310) );
  CMXI2X1 U22683 ( .A0(n12310), .A1(n12301), .S(n4080), .Z(n12317) );
  CMX2X1 U22684 ( .A0(n12302), .A1(n12317), .S(n3812), .Z(n12330) );
  CMXI2X1 U22685 ( .A0(n12303), .A1(n12330), .S(n3275), .Z(N6047) );
  CMX2X1 U22686 ( .A0(n12305), .A1(n12304), .S(n4315), .Z(n12567) );
  CMXI2X1 U22687 ( .A0(n12306), .A1(n12567), .S(n3438), .Z(N5246) );
  CMX2X1 U22688 ( .A0(N7375), .A1(N7374), .S(n3865), .Z(n12313) );
  CMXI2X1 U22689 ( .A0(n12313), .A1(n12307), .S(n4080), .Z(n12320) );
  CMX2X1 U22690 ( .A0(n12308), .A1(n12320), .S(n3771), .Z(n12333) );
  CMXI2X1 U22691 ( .A0(n12309), .A1(n12333), .S(n3438), .Z(N6048) );
  CMX2X1 U22692 ( .A0(N7374), .A1(N7373), .S(n3866), .Z(n12316) );
  CMXI2X1 U22693 ( .A0(n12316), .A1(n12310), .S(n4080), .Z(n12323) );
  CMX2X1 U22694 ( .A0(n12311), .A1(n12323), .S(n3805), .Z(n12336) );
  CMXI2X1 U22695 ( .A0(n12312), .A1(n12336), .S(n3438), .Z(N6049) );
  CMX2X1 U22696 ( .A0(N7373), .A1(N7372), .S(n3867), .Z(n12319) );
  CMXI2X1 U22697 ( .A0(n12319), .A1(n12313), .S(n4080), .Z(n12326) );
  CMX2X1 U22698 ( .A0(n12314), .A1(n12326), .S(n3807), .Z(n12344) );
  CMXI2X1 U22699 ( .A0(n12315), .A1(n12344), .S(n3438), .Z(N6050) );
  CMX2X1 U22700 ( .A0(N7372), .A1(N7371), .S(n3864), .Z(n12322) );
  CMXI2X1 U22701 ( .A0(n12322), .A1(n12316), .S(n4080), .Z(n12329) );
  CMX2X1 U22702 ( .A0(n12317), .A1(n12329), .S(n3808), .Z(n12347) );
  CMXI2X1 U22703 ( .A0(n12318), .A1(n12347), .S(n3438), .Z(N6051) );
  CMX2X1 U22704 ( .A0(N7371), .A1(N7370), .S(n3865), .Z(n12325) );
  CMXI2X1 U22705 ( .A0(n12325), .A1(n12319), .S(n4080), .Z(n12332) );
  CMX2X1 U22706 ( .A0(n12320), .A1(n12332), .S(n3809), .Z(n12350) );
  CMXI2X1 U22707 ( .A0(n12321), .A1(n12350), .S(n3438), .Z(N6052) );
  CMX2X1 U22708 ( .A0(N7370), .A1(N7369), .S(n3866), .Z(n12328) );
  CMXI2X1 U22709 ( .A0(n12328), .A1(n12322), .S(n4080), .Z(n12335) );
  CMX2X1 U22710 ( .A0(n12323), .A1(n12335), .S(n3810), .Z(n12353) );
  CMXI2X1 U22711 ( .A0(n12324), .A1(n12353), .S(n3437), .Z(N6053) );
  CMX2X1 U22712 ( .A0(N7369), .A1(N7368), .S(n3867), .Z(n12331) );
  CMXI2X1 U22713 ( .A0(n12331), .A1(n12325), .S(n4080), .Z(n12343) );
  CMX2X1 U22714 ( .A0(n12326), .A1(n12343), .S(n3811), .Z(n12356) );
  CMXI2X1 U22715 ( .A0(n12327), .A1(n12356), .S(n3437), .Z(N6054) );
  CMX2X1 U22716 ( .A0(N7368), .A1(N7367), .S(n3876), .Z(n12334) );
  CMXI2X1 U22717 ( .A0(n12334), .A1(n12328), .S(n4080), .Z(n12346) );
  CMX2X1 U22718 ( .A0(n12329), .A1(n12346), .S(n3812), .Z(n12359) );
  CMXI2X1 U22719 ( .A0(n12330), .A1(n12359), .S(n3437), .Z(N6055) );
  CMX2X1 U22720 ( .A0(N7367), .A1(N7366), .S(n3864), .Z(n12342) );
  CMXI2X1 U22721 ( .A0(n12342), .A1(n12331), .S(n4079), .Z(n12349) );
  CMX2X1 U22722 ( .A0(n12332), .A1(n12349), .S(n4319), .Z(n12362) );
  CMXI2X1 U22723 ( .A0(n12333), .A1(n12362), .S(n3437), .Z(N6056) );
  CMX2X1 U22724 ( .A0(N7366), .A1(N7365), .S(n3865), .Z(n12345) );
  CMXI2X1 U22725 ( .A0(n12345), .A1(n12334), .S(n4079), .Z(n12352) );
  CMX2X1 U22726 ( .A0(n12335), .A1(n12352), .S(n3771), .Z(n12365) );
  CMXI2X1 U22727 ( .A0(n12336), .A1(n12365), .S(n3437), .Z(N6057) );
  CMX2X1 U22728 ( .A0(n12338), .A1(n12337), .S(n3772), .Z(n12599) );
  CMXI2X1 U22729 ( .A0(n12339), .A1(n12599), .S(n3437), .Z(N5247) );
  CMXI2X1 U22730 ( .A0(n12341), .A1(n12340), .S(n3437), .Z(N5166) );
  CMX2X1 U22731 ( .A0(N7365), .A1(N7364), .S(n3866), .Z(n12348) );
  CMXI2X1 U22732 ( .A0(n12348), .A1(n12342), .S(n4079), .Z(n12355) );
  CMX2X1 U22733 ( .A0(n12343), .A1(n12355), .S(n3773), .Z(n12368) );
  CMXI2X1 U22734 ( .A0(n12344), .A1(n12368), .S(n3437), .Z(N6058) );
  CMX2X1 U22735 ( .A0(N7364), .A1(N7363), .S(n3867), .Z(n12351) );
  CMXI2X1 U22736 ( .A0(n12351), .A1(n12345), .S(n4079), .Z(n12358) );
  CMX2X1 U22737 ( .A0(n12346), .A1(n12358), .S(n3774), .Z(n12371) );
  CMXI2X1 U22738 ( .A0(n12347), .A1(n12371), .S(n3437), .Z(N6059) );
  CMX2X1 U22739 ( .A0(N7363), .A1(N7362), .S(n3868), .Z(n12354) );
  CMXI2X1 U22740 ( .A0(n12354), .A1(n12348), .S(n4079), .Z(n12361) );
  CMX2X1 U22741 ( .A0(n12349), .A1(n12361), .S(n3775), .Z(n12377) );
  CMXI2X1 U22742 ( .A0(n12350), .A1(n12377), .S(n3437), .Z(N6060) );
  CMX2X1 U22743 ( .A0(N7362), .A1(N7361), .S(n3869), .Z(n12357) );
  CMXI2X1 U22744 ( .A0(n12357), .A1(n12351), .S(n4079), .Z(n12364) );
  CMX2X1 U22745 ( .A0(n12352), .A1(n12364), .S(n3776), .Z(n12380) );
  CMXI2X1 U22746 ( .A0(n12353), .A1(n12380), .S(n3436), .Z(N6061) );
  CMX2X1 U22747 ( .A0(N7361), .A1(N7360), .S(n3870), .Z(n12360) );
  CMXI2X1 U22748 ( .A0(n12360), .A1(n12354), .S(n4079), .Z(n12367) );
  CMX2X1 U22749 ( .A0(n12355), .A1(n12367), .S(n3777), .Z(n12383) );
  CMXI2X1 U22750 ( .A0(n12356), .A1(n12383), .S(n3436), .Z(N6062) );
  CMX2X1 U22751 ( .A0(N7360), .A1(N7359), .S(n3872), .Z(n12363) );
  CMXI2X1 U22752 ( .A0(n12363), .A1(n12357), .S(n4079), .Z(n12370) );
  CMX2X1 U22753 ( .A0(n12358), .A1(n12370), .S(n3790), .Z(n12386) );
  CMX2X1 U22754 ( .A0(N7359), .A1(N7358), .S(n3873), .Z(n12366) );
  CMXI2X1 U22755 ( .A0(n12366), .A1(n12360), .S(n4079), .Z(n12376) );
  CMX2X1 U22756 ( .A0(n12361), .A1(n12376), .S(n3791), .Z(n12389) );
  CMX2X1 U22757 ( .A0(N7358), .A1(N7357), .S(n3871), .Z(n12369) );
  CMXI2X1 U22758 ( .A0(n12369), .A1(n12363), .S(n4079), .Z(n12379) );
  CMX2X1 U22759 ( .A0(n12364), .A1(n12379), .S(n3773), .Z(n12392) );
  CMXI2X1 U22760 ( .A0(n12365), .A1(n12392), .S(n3439), .Z(N6065) );
  CMX2X1 U22761 ( .A0(N7357), .A1(N7356), .S(n3872), .Z(n12375) );
  CMXI2X1 U22762 ( .A0(n12375), .A1(n12366), .S(n4079), .Z(n12382) );
  CMX2X1 U22763 ( .A0(n12367), .A1(n12382), .S(n3774), .Z(n12395) );
  CMXI2X1 U22764 ( .A0(n12368), .A1(n12395), .S(n3439), .Z(N6066) );
  CMX2X1 U22765 ( .A0(N7356), .A1(N7355), .S(n3868), .Z(n12378) );
  CMXI2X1 U22766 ( .A0(n12378), .A1(n12369), .S(n4079), .Z(n12385) );
  CMX2X1 U22767 ( .A0(n12370), .A1(n12385), .S(n3772), .Z(n12398) );
  CMXI2X1 U22768 ( .A0(n12371), .A1(n12398), .S(n3439), .Z(N6067) );
  CMX2X1 U22769 ( .A0(n12373), .A1(n12372), .S(n3773), .Z(n12633) );
  CMXI2X1 U22770 ( .A0(n12374), .A1(n12633), .S(n3439), .Z(N5248) );
  CMX2X1 U22771 ( .A0(N7355), .A1(N7354), .S(n3869), .Z(n12381) );
  CMXI2X1 U22772 ( .A0(n12381), .A1(n12375), .S(n4079), .Z(n12388) );
  CMX2X1 U22773 ( .A0(n12376), .A1(n12388), .S(n3774), .Z(n12401) );
  CMXI2X1 U22774 ( .A0(n12377), .A1(n12401), .S(n3439), .Z(N6068) );
  CMX2X1 U22775 ( .A0(N7354), .A1(N7353), .S(n3870), .Z(n12384) );
  CMXI2X1 U22776 ( .A0(n12384), .A1(n12378), .S(n4079), .Z(n12391) );
  CMX2X1 U22777 ( .A0(n12379), .A1(n12391), .S(n3775), .Z(n12404) );
  CMXI2X1 U22778 ( .A0(n12380), .A1(n12404), .S(n3439), .Z(N6069) );
  CMX2X1 U22779 ( .A0(N7353), .A1(N7352), .S(n3871), .Z(n12387) );
  CMXI2X1 U22780 ( .A0(n12387), .A1(n12381), .S(n4079), .Z(n12394) );
  CMX2X1 U22781 ( .A0(n12382), .A1(n12394), .S(n3776), .Z(n12410) );
  CMXI2X1 U22782 ( .A0(n12383), .A1(n12410), .S(n3439), .Z(N6070) );
  CMX2X1 U22783 ( .A0(N7352), .A1(N7351), .S(n3868), .Z(n12390) );
  CMXI2X1 U22784 ( .A0(n12390), .A1(n12384), .S(n4079), .Z(n12397) );
  CMX2X1 U22785 ( .A0(n12385), .A1(n12397), .S(n3806), .Z(n12413) );
  CMXI2X1 U22786 ( .A0(n12386), .A1(n12413), .S(n3439), .Z(N6071) );
  CMX2X1 U22787 ( .A0(N7351), .A1(N7350), .S(n3869), .Z(n12393) );
  CMXI2X1 U22788 ( .A0(n12393), .A1(n12387), .S(n4078), .Z(n12400) );
  CMX2X1 U22789 ( .A0(n12388), .A1(n12400), .S(n3791), .Z(n12416) );
  CMX2X1 U22790 ( .A0(N7350), .A1(N7349), .S(n3870), .Z(n12396) );
  CMXI2X1 U22791 ( .A0(n12396), .A1(n12390), .S(n4078), .Z(n12403) );
  CMX2X1 U22792 ( .A0(n12391), .A1(n12403), .S(n3792), .Z(n12419) );
  CMXI2X1 U22793 ( .A0(n12392), .A1(n12419), .S(n3439), .Z(N6073) );
  CMX2X1 U22794 ( .A0(N7349), .A1(N7348), .S(n3871), .Z(n12399) );
  CMXI2X1 U22795 ( .A0(n12399), .A1(n12393), .S(n4078), .Z(n12409) );
  CMX2X1 U22796 ( .A0(n12394), .A1(n12409), .S(n3793), .Z(n12422) );
  CMXI2X1 U22797 ( .A0(n12395), .A1(n12422), .S(n3439), .Z(N6074) );
  CMX2X1 U22798 ( .A0(N7348), .A1(N7347), .S(n3877), .Z(n12402) );
  CMXI2X1 U22799 ( .A0(n12402), .A1(n12396), .S(n4078), .Z(n12412) );
  CMX2X1 U22800 ( .A0(n12397), .A1(n12412), .S(n3794), .Z(n12425) );
  CMXI2X1 U22801 ( .A0(n12398), .A1(n12425), .S(n3438), .Z(N6075) );
  CMX2X1 U22802 ( .A0(N7347), .A1(N7346), .S(n3873), .Z(n12408) );
  CMXI2X1 U22803 ( .A0(n12408), .A1(n12399), .S(n4078), .Z(n12415) );
  CMX2X1 U22804 ( .A0(n12400), .A1(n12415), .S(n3795), .Z(n12428) );
  CMXI2X1 U22805 ( .A0(n12401), .A1(n12428), .S(n3438), .Z(N6076) );
  CMX2X1 U22806 ( .A0(N7346), .A1(N7345), .S(n3874), .Z(n12411) );
  CMXI2X1 U22807 ( .A0(n12411), .A1(n12402), .S(n4078), .Z(n12418) );
  CMX2X1 U22808 ( .A0(n12403), .A1(n12418), .S(n3796), .Z(n12431) );
  CMXI2X1 U22809 ( .A0(n12404), .A1(n12431), .S(n3438), .Z(N6077) );
  CMX2X1 U22810 ( .A0(n12406), .A1(n12405), .S(n3797), .Z(n12657) );
  CMXI2X1 U22811 ( .A0(n12407), .A1(n12657), .S(n3438), .Z(N5249) );
  CMX2X1 U22812 ( .A0(N7345), .A1(N7344), .S(n3875), .Z(n12414) );
  CMXI2X1 U22813 ( .A0(n12414), .A1(n12408), .S(n4078), .Z(n12421) );
  CMX2X1 U22814 ( .A0(n12409), .A1(n12421), .S(n3805), .Z(n12434) );
  CMXI2X1 U22815 ( .A0(n12410), .A1(n12434), .S(n3438), .Z(N6078) );
  CMX2X1 U22816 ( .A0(N7344), .A1(N7343), .S(n3876), .Z(n12417) );
  CMXI2X1 U22817 ( .A0(n12417), .A1(n12411), .S(n4078), .Z(n12424) );
  CMX2X1 U22818 ( .A0(n12412), .A1(n12424), .S(n3806), .Z(n12437) );
  CMXI2X1 U22819 ( .A0(n12413), .A1(n12437), .S(n3441), .Z(N6079) );
  CMX2X1 U22820 ( .A0(N7343), .A1(N7342), .S(n3877), .Z(n12420) );
  CMXI2X1 U22821 ( .A0(n12420), .A1(n12414), .S(n4078), .Z(n12427) );
  CMX2X1 U22822 ( .A0(n12415), .A1(n12427), .S(n3773), .Z(n12442) );
  CMXI2X1 U22823 ( .A0(n12416), .A1(n12442), .S(n3441), .Z(N6080) );
  CMX2X1 U22824 ( .A0(N7342), .A1(N7341), .S(n3878), .Z(n12423) );
  CMXI2X1 U22825 ( .A0(n12423), .A1(n12417), .S(n4078), .Z(n12430) );
  CMX2X1 U22826 ( .A0(n12418), .A1(n12430), .S(n3809), .Z(n12445) );
  CMXI2X1 U22827 ( .A0(n12419), .A1(n12445), .S(n3441), .Z(N6081) );
  CMX2X1 U22828 ( .A0(N7341), .A1(N7340), .S(n3879), .Z(n12426) );
  CMXI2X1 U22829 ( .A0(n12426), .A1(n12420), .S(n4078), .Z(n12433) );
  CMX2X1 U22830 ( .A0(n12421), .A1(n12433), .S(n3809), .Z(n12448) );
  CMXI2X1 U22831 ( .A0(n12422), .A1(n12448), .S(n3441), .Z(N6082) );
  CMX2X1 U22832 ( .A0(N7340), .A1(N7339), .S(n3874), .Z(n12429) );
  CMXI2X1 U22833 ( .A0(n12429), .A1(n12423), .S(n4078), .Z(n12436) );
  CMX2X1 U22834 ( .A0(n12424), .A1(n12436), .S(n3810), .Z(n12451) );
  CMXI2X1 U22835 ( .A0(n12425), .A1(n12451), .S(n3441), .Z(N6083) );
  CMX2X1 U22836 ( .A0(N7339), .A1(N7338), .S(n3875), .Z(n12432) );
  CMXI2X1 U22837 ( .A0(n12432), .A1(n12426), .S(n4078), .Z(n12441) );
  CMX2X1 U22838 ( .A0(n12427), .A1(n12441), .S(n3811), .Z(n12454) );
  CMXI2X1 U22839 ( .A0(n12428), .A1(n12454), .S(n3441), .Z(N6084) );
  CMX2X1 U22840 ( .A0(N7338), .A1(N7337), .S(n3880), .Z(n12435) );
  CMXI2X1 U22841 ( .A0(n12435), .A1(n12429), .S(n4078), .Z(n12444) );
  CMX2X1 U22842 ( .A0(n12430), .A1(n12444), .S(n3812), .Z(n12457) );
  CMXI2X1 U22843 ( .A0(n12431), .A1(n12457), .S(n3441), .Z(N6085) );
  CMX2X1 U22844 ( .A0(N7337), .A1(N7336), .S(n3881), .Z(n12440) );
  CMXI2X1 U22845 ( .A0(n12440), .A1(n12432), .S(n4078), .Z(n12447) );
  CMX2X1 U22846 ( .A0(n12433), .A1(n12447), .S(n4308), .Z(n12460) );
  CMXI2X1 U22847 ( .A0(n12434), .A1(n12460), .S(n3441), .Z(N6086) );
  CMX2X1 U22848 ( .A0(N7336), .A1(N7335), .S(n3872), .Z(n12443) );
  CMXI2X1 U22849 ( .A0(n12443), .A1(n12435), .S(n4078), .Z(n12450) );
  CMX2X1 U22850 ( .A0(n12436), .A1(n12450), .S(n3809), .Z(n12463) );
  CMXI2X1 U22851 ( .A0(n12437), .A1(n12463), .S(n3441), .Z(N6087) );
  CMXI2X1 U22852 ( .A0(n12439), .A1(n12438), .S(n3440), .Z(N5250) );
  CMX2X1 U22853 ( .A0(N7335), .A1(N7334), .S(n3873), .Z(n12446) );
  CMXI2X1 U22854 ( .A0(n12446), .A1(n12440), .S(n4077), .Z(n12453) );
  CMX2X1 U22855 ( .A0(n12441), .A1(n12453), .S(n3807), .Z(n12466) );
  CMXI2X1 U22856 ( .A0(n12442), .A1(n12466), .S(n3440), .Z(N6088) );
  CMX2X1 U22857 ( .A0(N7334), .A1(N7333), .S(n3874), .Z(n12449) );
  CMXI2X1 U22858 ( .A0(n12449), .A1(n12443), .S(n4077), .Z(n12456) );
  CMX2X1 U22859 ( .A0(n12444), .A1(n12456), .S(n3808), .Z(n12469) );
  CMXI2X1 U22860 ( .A0(n12445), .A1(n12469), .S(n3440), .Z(N6089) );
  CMX2X1 U22861 ( .A0(N7333), .A1(N7332), .S(n3875), .Z(n12452) );
  CMXI2X1 U22862 ( .A0(n12452), .A1(n12446), .S(n4077), .Z(n12459) );
  CMX2X1 U22863 ( .A0(n12447), .A1(n12459), .S(n3809), .Z(n12474) );
  CMXI2X1 U22864 ( .A0(n12448), .A1(n12474), .S(n3440), .Z(N6090) );
  CMX2X1 U22865 ( .A0(N7332), .A1(N7331), .S(n3872), .Z(n12455) );
  CMXI2X1 U22866 ( .A0(n12455), .A1(n12449), .S(n4077), .Z(n12462) );
  CMX2X1 U22867 ( .A0(n12450), .A1(n12462), .S(n3810), .Z(n12477) );
  CMXI2X1 U22868 ( .A0(n12451), .A1(n12477), .S(n3440), .Z(N6091) );
  CMX2X1 U22869 ( .A0(N7331), .A1(N7330), .S(n3873), .Z(n12458) );
  CMXI2X1 U22870 ( .A0(n12458), .A1(n12452), .S(n4077), .Z(n12465) );
  CMX2X1 U22871 ( .A0(n12453), .A1(n12465), .S(n3811), .Z(n12480) );
  CMXI2X1 U22872 ( .A0(n12454), .A1(n12480), .S(n3440), .Z(N6092) );
  CMX2X1 U22873 ( .A0(N7330), .A1(N7329), .S(n3874), .Z(n12461) );
  CMXI2X1 U22874 ( .A0(n12461), .A1(n12455), .S(n4077), .Z(n12468) );
  CMX2X1 U22875 ( .A0(n12456), .A1(n12468), .S(n3806), .Z(n12483) );
  CMXI2X1 U22876 ( .A0(n12457), .A1(n12483), .S(n3440), .Z(N6093) );
  CMX2X1 U22877 ( .A0(N7329), .A1(N7328), .S(n3875), .Z(n12464) );
  CMXI2X1 U22878 ( .A0(n12464), .A1(n12458), .S(n4077), .Z(n12473) );
  CMX2X1 U22879 ( .A0(n12459), .A1(n12473), .S(n3812), .Z(n12486) );
  CMXI2X1 U22880 ( .A0(n12460), .A1(n12486), .S(n3440), .Z(N6094) );
  CMX2X1 U22881 ( .A0(N7328), .A1(N7327), .S(n3878), .Z(n12467) );
  CMXI2X1 U22882 ( .A0(n12467), .A1(n12461), .S(n4077), .Z(n12476) );
  CMX2X1 U22883 ( .A0(n12462), .A1(n12476), .S(n4308), .Z(n12489) );
  CMXI2X1 U22884 ( .A0(n12463), .A1(n12489), .S(n3440), .Z(N6095) );
  CMX2X1 U22885 ( .A0(N7327), .A1(N7326), .S(n3862), .Z(n12472) );
  CMXI2X1 U22886 ( .A0(n12472), .A1(n12464), .S(n4077), .Z(n12479) );
  CMX2X1 U22887 ( .A0(n12465), .A1(n12479), .S(n3776), .Z(n12492) );
  CMXI2X1 U22888 ( .A0(n12466), .A1(n12492), .S(n3443), .Z(N6096) );
  CMX2X1 U22889 ( .A0(N7326), .A1(N7325), .S(n3863), .Z(n12475) );
  CMXI2X1 U22890 ( .A0(n12475), .A1(n12467), .S(n4077), .Z(n12482) );
  CMX2X1 U22891 ( .A0(n12468), .A1(n12482), .S(n3777), .Z(n12495) );
  CMXI2X1 U22892 ( .A0(n12469), .A1(n12495), .S(n3443), .Z(N6097) );
  CMXI2X1 U22893 ( .A0(n12471), .A1(n12470), .S(n3443), .Z(N5251) );
  CMX2X1 U22894 ( .A0(N7325), .A1(N7324), .S(n3864), .Z(n12478) );
  CMXI2X1 U22895 ( .A0(n12478), .A1(n12472), .S(n4077), .Z(n12485) );
  CMX2X1 U22896 ( .A0(n12473), .A1(n12485), .S(n3790), .Z(n12498) );
  CMXI2X1 U22897 ( .A0(n12474), .A1(n12498), .S(n3443), .Z(N6098) );
  CMX2X1 U22898 ( .A0(N7324), .A1(N7323), .S(n3865), .Z(n12481) );
  CMXI2X1 U22899 ( .A0(n12481), .A1(n12475), .S(n4077), .Z(n12488) );
  CMX2X1 U22900 ( .A0(n12476), .A1(n12488), .S(n3791), .Z(n12501) );
  CMXI2X1 U22901 ( .A0(n12477), .A1(n12501), .S(n3443), .Z(N6099) );
  CMX2X1 U22902 ( .A0(N7323), .A1(N7322), .S(n3866), .Z(n12484) );
  CMXI2X1 U22903 ( .A0(n12484), .A1(n12478), .S(n4077), .Z(n12491) );
  CMX2X1 U22904 ( .A0(n12479), .A1(n12491), .S(n3792), .Z(n12506) );
  CMXI2X1 U22905 ( .A0(n12480), .A1(n12506), .S(n3442), .Z(N6100) );
  CMX2X1 U22906 ( .A0(N7322), .A1(N7321), .S(n3867), .Z(n12487) );
  CMXI2X1 U22907 ( .A0(n12487), .A1(n12481), .S(n4077), .Z(n12494) );
  CMX2X1 U22908 ( .A0(n12482), .A1(n12494), .S(n3795), .Z(n12509) );
  CMXI2X1 U22909 ( .A0(n12483), .A1(n12509), .S(n3442), .Z(N6101) );
  CMX2X1 U22910 ( .A0(N7321), .A1(N7320), .S(n3868), .Z(n12490) );
  CMXI2X1 U22911 ( .A0(n12490), .A1(n12484), .S(n4077), .Z(n12497) );
  CMX2X1 U22912 ( .A0(n12485), .A1(n12497), .S(n3807), .Z(n12512) );
  CMXI2X1 U22913 ( .A0(n12486), .A1(n12512), .S(n3442), .Z(N6102) );
  CMX2X1 U22914 ( .A0(N7320), .A1(N7319), .S(n3876), .Z(n12493) );
  CMXI2X1 U22915 ( .A0(n12493), .A1(n12487), .S(n4077), .Z(n12500) );
  CMX2X1 U22916 ( .A0(n12488), .A1(n12500), .S(n3808), .Z(n12515) );
  CMXI2X1 U22917 ( .A0(n12489), .A1(n12515), .S(n3442), .Z(N6103) );
  CMX2X1 U22918 ( .A0(N7319), .A1(N7318), .S(n3877), .Z(n12496) );
  CMXI2X1 U22919 ( .A0(n12496), .A1(n12490), .S(n4076), .Z(n12505) );
  CMX2X1 U22920 ( .A0(n12491), .A1(n12505), .S(n3809), .Z(n12518) );
  CMXI2X1 U22921 ( .A0(n12492), .A1(n12518), .S(n3442), .Z(N6104) );
  CMX2X1 U22922 ( .A0(N7318), .A1(N7317), .S(n3869), .Z(n12499) );
  CMXI2X1 U22923 ( .A0(n12499), .A1(n12493), .S(n4076), .Z(n12508) );
  CMX2X1 U22924 ( .A0(n12494), .A1(n12508), .S(n3810), .Z(n12521) );
  CMXI2X1 U22925 ( .A0(n12495), .A1(n12521), .S(n3442), .Z(N6105) );
  CMX2X1 U22926 ( .A0(N7317), .A1(N7316), .S(n3870), .Z(n12504) );
  CMXI2X1 U22927 ( .A0(n12504), .A1(n12496), .S(n4076), .Z(n12511) );
  CMX2X1 U22928 ( .A0(n12497), .A1(n12511), .S(n3811), .Z(n12524) );
  CMXI2X1 U22929 ( .A0(n12498), .A1(n12524), .S(n3442), .Z(N6106) );
  CMX2X1 U22930 ( .A0(N7316), .A1(N7315), .S(n3876), .Z(n12507) );
  CMXI2X1 U22931 ( .A0(n12507), .A1(n12499), .S(n4076), .Z(n12514) );
  CMX2X1 U22932 ( .A0(n12500), .A1(n12514), .S(n3812), .Z(n12527) );
  CMXI2X1 U22933 ( .A0(n12501), .A1(n12527), .S(n3442), .Z(N6107) );
  CMXI2X1 U22934 ( .A0(n12503), .A1(n12502), .S(n3442), .Z(N5252) );
  CMX2X1 U22935 ( .A0(N7315), .A1(N7314), .S(n3877), .Z(n12510) );
  CMXI2X1 U22936 ( .A0(n12510), .A1(n12504), .S(n4076), .Z(n12517) );
  CMX2X1 U22937 ( .A0(n12505), .A1(n12517), .S(n4323), .Z(n12530) );
  CMXI2X1 U22938 ( .A0(n12506), .A1(n12530), .S(n3442), .Z(N6108) );
  CMX2X1 U22939 ( .A0(N7314), .A1(N7313), .S(n3878), .Z(n12513) );
  CMXI2X1 U22940 ( .A0(n12513), .A1(n12507), .S(n4076), .Z(n12520) );
  CMX2X1 U22941 ( .A0(n12508), .A1(n12520), .S(n3771), .Z(n12533) );
  CMXI2X1 U22942 ( .A0(n12509), .A1(n12533), .S(n3442), .Z(N6109) );
  CMX2X1 U22943 ( .A0(N7313), .A1(N7312), .S(n3879), .Z(n12516) );
  CMXI2X1 U22944 ( .A0(n12516), .A1(n12510), .S(n4076), .Z(n12523) );
  CMX2X1 U22945 ( .A0(n12511), .A1(n12523), .S(n3772), .Z(n12538) );
  CMXI2X1 U22946 ( .A0(n12512), .A1(n12538), .S(n3441), .Z(N6110) );
  CMX2X1 U22947 ( .A0(N7312), .A1(N7311), .S(n3876), .Z(n12519) );
  CMXI2X1 U22948 ( .A0(n12519), .A1(n12513), .S(n4076), .Z(n12526) );
  CMX2X1 U22949 ( .A0(n12514), .A1(n12526), .S(n3773), .Z(n12541) );
  CMXI2X1 U22950 ( .A0(n12515), .A1(n12541), .S(n3441), .Z(N6111) );
  CMX2X1 U22951 ( .A0(N7311), .A1(N7310), .S(n3877), .Z(n12522) );
  CMXI2X1 U22952 ( .A0(n12522), .A1(n12516), .S(n4076), .Z(n12529) );
  CMX2X1 U22953 ( .A0(n12517), .A1(n12529), .S(n3774), .Z(n12544) );
  CMXI2X1 U22954 ( .A0(n12518), .A1(n12544), .S(n3445), .Z(N6112) );
  CMX2X1 U22955 ( .A0(N7310), .A1(N7309), .S(n3878), .Z(n12525) );
  CMXI2X1 U22956 ( .A0(n12525), .A1(n12519), .S(n4076), .Z(n12532) );
  CMX2X1 U22957 ( .A0(n12520), .A1(n12532), .S(n3775), .Z(n12547) );
  CMXI2X1 U22958 ( .A0(n12521), .A1(n12547), .S(n3444), .Z(N6113) );
  CMX2X1 U22959 ( .A0(N7309), .A1(N7308), .S(n3879), .Z(n12528) );
  CMXI2X1 U22960 ( .A0(n12528), .A1(n12522), .S(n4076), .Z(n12537) );
  CMX2X1 U22961 ( .A0(n12523), .A1(n12537), .S(n3776), .Z(n12550) );
  CMXI2X1 U22962 ( .A0(n12524), .A1(n12550), .S(n3444), .Z(N6114) );
  CMX2X1 U22963 ( .A0(N7308), .A1(N7307), .S(n3879), .Z(n12531) );
  CMXI2X1 U22964 ( .A0(n12531), .A1(n12525), .S(n4076), .Z(n12540) );
  CMX2X1 U22965 ( .A0(n12526), .A1(n12540), .S(n3777), .Z(n12553) );
  CMXI2X1 U22966 ( .A0(n12527), .A1(n12553), .S(n3444), .Z(N6115) );
  CMX2X1 U22967 ( .A0(N7307), .A1(N7306), .S(n3871), .Z(n12536) );
  CMXI2X1 U22968 ( .A0(n12536), .A1(n12528), .S(n4076), .Z(n12543) );
  CMX2X1 U22969 ( .A0(n12529), .A1(n12543), .S(n3790), .Z(n12556) );
  CMXI2X1 U22970 ( .A0(n12530), .A1(n12556), .S(n3444), .Z(N6116) );
  CMX2X1 U22971 ( .A0(N7306), .A1(N7305), .S(n3872), .Z(n12539) );
  CMXI2X1 U22972 ( .A0(n12539), .A1(n12531), .S(n4076), .Z(n12546) );
  CMX2X1 U22973 ( .A0(n12532), .A1(n12546), .S(n3791), .Z(n12559) );
  CMXI2X1 U22974 ( .A0(n12533), .A1(n12559), .S(n3444), .Z(N6117) );
  CMXI2X1 U22975 ( .A0(n12535), .A1(n12534), .S(n3444), .Z(N5253) );
  CMX2X1 U22976 ( .A0(N7305), .A1(N7304), .S(n3873), .Z(n12542) );
  CMXI2X1 U22977 ( .A0(n12542), .A1(n12536), .S(n4076), .Z(n12549) );
  CMX2X1 U22978 ( .A0(n12537), .A1(n12549), .S(n4310), .Z(n12562) );
  CMXI2X1 U22979 ( .A0(n12538), .A1(n12562), .S(n3444), .Z(N6118) );
  CMX2X1 U22980 ( .A0(N7304), .A1(N7303), .S(n3874), .Z(n12545) );
  CMXI2X1 U22981 ( .A0(n12545), .A1(n12539), .S(n4076), .Z(n12552) );
  CMX2X1 U22982 ( .A0(n12540), .A1(n12552), .S(n3771), .Z(n12565) );
  CMXI2X1 U22983 ( .A0(n12541), .A1(n12565), .S(n3444), .Z(N6119) );
  CMX2X1 U22984 ( .A0(N7303), .A1(N7302), .S(n3875), .Z(n12548) );
  CMXI2X1 U22985 ( .A0(n12548), .A1(n12542), .S(n4075), .Z(n12555) );
  CMX2X1 U22986 ( .A0(n12543), .A1(n12555), .S(n3793), .Z(n12570) );
  CMXI2X1 U22987 ( .A0(n12544), .A1(n12570), .S(n3444), .Z(N6120) );
  CMX2X1 U22988 ( .A0(N7302), .A1(N7301), .S(n3876), .Z(n12551) );
  CMXI2X1 U22989 ( .A0(n12551), .A1(n12545), .S(n4075), .Z(n12558) );
  CMX2X1 U22990 ( .A0(n12546), .A1(n12558), .S(n3794), .Z(n12573) );
  CMXI2X1 U22991 ( .A0(n12547), .A1(n12573), .S(n3444), .Z(N6121) );
  CMX2X1 U22992 ( .A0(N7301), .A1(N7300), .S(n3877), .Z(n12554) );
  CMXI2X1 U22993 ( .A0(n12554), .A1(n12548), .S(n4075), .Z(n12561) );
  CMX2X1 U22994 ( .A0(n12549), .A1(n12561), .S(n3795), .Z(n12576) );
  CMXI2X1 U22995 ( .A0(n12550), .A1(n12576), .S(n3444), .Z(N6122) );
  CMX2X1 U22996 ( .A0(N7300), .A1(N7299), .S(n3868), .Z(n12557) );
  CMXI2X1 U22997 ( .A0(n12557), .A1(n12551), .S(n4075), .Z(n12564) );
  CMX2X1 U22998 ( .A0(n12552), .A1(n12564), .S(n3796), .Z(n12579) );
  CMXI2X1 U22999 ( .A0(n12553), .A1(n12579), .S(n3443), .Z(N6123) );
  CMX2X1 U23000 ( .A0(N7299), .A1(N7298), .S(n3866), .Z(n12560) );
  CMXI2X1 U23001 ( .A0(n12560), .A1(n12554), .S(n4075), .Z(n12569) );
  CMX2X1 U23002 ( .A0(n12555), .A1(n12569), .S(n3797), .Z(n12582) );
  CMXI2X1 U23003 ( .A0(n12556), .A1(n12582), .S(n3443), .Z(N6124) );
  CMX2X1 U23004 ( .A0(N7298), .A1(N7297), .S(n3867), .Z(n12563) );
  CMXI2X1 U23005 ( .A0(n12563), .A1(n12557), .S(n4075), .Z(n12572) );
  CMX2X1 U23006 ( .A0(n12558), .A1(n12572), .S(n3796), .Z(n12585) );
  CMXI2X1 U23007 ( .A0(n12559), .A1(n12585), .S(n3443), .Z(N6125) );
  CMX2X1 U23008 ( .A0(N7297), .A1(N7296), .S(n3869), .Z(n12568) );
  CMXI2X1 U23009 ( .A0(n12568), .A1(n12560), .S(n4075), .Z(n12575) );
  CMX2X1 U23010 ( .A0(n12561), .A1(n12575), .S(n3792), .Z(n12588) );
  CMXI2X1 U23011 ( .A0(n12562), .A1(n12588), .S(n3443), .Z(N6126) );
  CMX2X1 U23012 ( .A0(N7296), .A1(N7295), .S(n3870), .Z(n12571) );
  CMXI2X1 U23013 ( .A0(n12571), .A1(n12563), .S(n4075), .Z(n12578) );
  CMX2X1 U23014 ( .A0(n12564), .A1(n12578), .S(n3793), .Z(n12591) );
  CMXI2X1 U23015 ( .A0(n12565), .A1(n12591), .S(n3443), .Z(N6127) );
  CMXI2X1 U23016 ( .A0(n12567), .A1(n12566), .S(n3424), .Z(N5254) );
  CMX2X1 U23017 ( .A0(N7295), .A1(N7294), .S(n3862), .Z(n12574) );
  CMXI2X1 U23018 ( .A0(n12574), .A1(n12568), .S(n4075), .Z(n12581) );
  CMX2X1 U23019 ( .A0(n12569), .A1(n12581), .S(n3794), .Z(n12594) );
  CMXI2X1 U23020 ( .A0(n12570), .A1(n12594), .S(n3463), .Z(N6128) );
  CMX2X1 U23021 ( .A0(N7294), .A1(N7293), .S(n3863), .Z(n12577) );
  CMXI2X1 U23022 ( .A0(n12577), .A1(n12571), .S(n4075), .Z(n12584) );
  CMX2X1 U23023 ( .A0(n12572), .A1(n12584), .S(n3795), .Z(n12597) );
  CMXI2X1 U23024 ( .A0(n12573), .A1(n12597), .S(n3446), .Z(N6129) );
  CMX2X1 U23025 ( .A0(N7293), .A1(N7292), .S(n3864), .Z(n12580) );
  CMXI2X1 U23026 ( .A0(n12580), .A1(n12574), .S(n4075), .Z(n12587) );
  CMX2X1 U23027 ( .A0(n12575), .A1(n12587), .S(n3796), .Z(n12602) );
  CMXI2X1 U23028 ( .A0(n12576), .A1(n12602), .S(n3446), .Z(N6130) );
  CMX2X1 U23029 ( .A0(N7292), .A1(N7291), .S(n3865), .Z(n12583) );
  CMXI2X1 U23030 ( .A0(n12583), .A1(n12577), .S(n4075), .Z(n12590) );
  CMX2X1 U23031 ( .A0(n12578), .A1(n12590), .S(n3797), .Z(n12605) );
  CMXI2X1 U23032 ( .A0(n12579), .A1(n12605), .S(n3446), .Z(N6131) );
  CMX2X1 U23033 ( .A0(N7291), .A1(N7290), .S(n3878), .Z(n12586) );
  CMXI2X1 U23034 ( .A0(n12586), .A1(n12580), .S(n4075), .Z(n12593) );
  CMX2X1 U23035 ( .A0(n12581), .A1(n12593), .S(n3805), .Z(n12608) );
  CMXI2X1 U23036 ( .A0(n12582), .A1(n12608), .S(n3446), .Z(N6132) );
  CMX2X1 U23037 ( .A0(N7290), .A1(N7289), .S(n3879), .Z(n12589) );
  CMXI2X1 U23038 ( .A0(n12589), .A1(n12583), .S(n4075), .Z(n12596) );
  CMX2X1 U23039 ( .A0(n12584), .A1(n12596), .S(n3806), .Z(n12611) );
  CMXI2X1 U23040 ( .A0(n12585), .A1(n12611), .S(n3446), .Z(N6133) );
  CMX2X1 U23041 ( .A0(N7289), .A1(N7288), .S(n3880), .Z(n12592) );
  CMXI2X1 U23042 ( .A0(n12592), .A1(n12586), .S(n4075), .Z(n12601) );
  CMX2X1 U23043 ( .A0(n12587), .A1(n12601), .S(n3807), .Z(n12614) );
  CMXI2X1 U23044 ( .A0(n12588), .A1(n12614), .S(n3446), .Z(N6134) );
  CMX2X1 U23045 ( .A0(N7288), .A1(N7287), .S(n3881), .Z(n12595) );
  CMXI2X1 U23046 ( .A0(n12595), .A1(n12589), .S(n4075), .Z(n12604) );
  CMX2X1 U23047 ( .A0(n12590), .A1(n12604), .S(n3808), .Z(n12617) );
  CMXI2X1 U23048 ( .A0(n12591), .A1(n12617), .S(n3445), .Z(N6135) );
  CMXI2X1 U23049 ( .A0(n12600), .A1(n12592), .S(n4074), .Z(n12607) );
  CMX2X1 U23050 ( .A0(n12593), .A1(n12607), .S(n3809), .Z(n12621) );
  CMXI2X1 U23051 ( .A0(n12594), .A1(n12621), .S(n3445), .Z(N6136) );
  CMXI2X1 U23052 ( .A0(n12603), .A1(n12595), .S(n4074), .Z(n12610) );
  CMX2X1 U23053 ( .A0(n12596), .A1(n12610), .S(n3810), .Z(n12625) );
  CMXI2X1 U23054 ( .A0(n12597), .A1(n12625), .S(n3445), .Z(N6137) );
  CMXI2X1 U23055 ( .A0(n12599), .A1(n12598), .S(n3445), .Z(N5255) );
  CMXI2X1 U23056 ( .A0(n12606), .A1(n12600), .S(n4074), .Z(n12613) );
  CMX2X1 U23057 ( .A0(n12601), .A1(n12613), .S(n3811), .Z(n12628) );
  CMXI2X1 U23058 ( .A0(n12602), .A1(n12628), .S(n3445), .Z(N6138) );
  CMXI2X1 U23059 ( .A0(n12609), .A1(n12603), .S(n4074), .Z(n12616) );
  CMX2X1 U23060 ( .A0(n12604), .A1(n12616), .S(n3812), .Z(n12631) );
  CMXI2X1 U23061 ( .A0(n12605), .A1(n12631), .S(n3445), .Z(N6139) );
  CMXI2X1 U23062 ( .A0(n12612), .A1(n12606), .S(n4074), .Z(n12620) );
  CMX2X1 U23063 ( .A0(n12607), .A1(n12620), .S(n4321), .Z(n12636) );
  CMXI2X1 U23064 ( .A0(n12608), .A1(n12636), .S(n3445), .Z(N6140) );
  CMXI2X1 U23065 ( .A0(n12615), .A1(n12609), .S(n4074), .Z(n12624) );
  CMX2X1 U23066 ( .A0(n12610), .A1(n12624), .S(n3771), .Z(n12639) );
  CMXI2X1 U23067 ( .A0(n12611), .A1(n12639), .S(n3445), .Z(N6141) );
  CMXI2X1 U23068 ( .A0(n12618), .A1(n12612), .S(n4074), .Z(n12627) );
  CMX2X1 U23069 ( .A0(n12613), .A1(n12627), .S(n3771), .Z(n12641) );
  CMXI2X1 U23070 ( .A0(n12614), .A1(n12641), .S(n3445), .Z(N6142) );
  CMXI2X1 U23071 ( .A0(n12622), .A1(n12615), .S(n4074), .Z(n12630) );
  CMX2X1 U23072 ( .A0(n12616), .A1(n12630), .S(n3772), .Z(n12643) );
  CMXI2X1 U23073 ( .A0(n12619), .A1(n12618), .S(n4074), .Z(n12635) );
  CMX2X1 U23074 ( .A0(n12620), .A1(n12635), .S(n3805), .Z(n12645) );
  CMXI2X1 U23075 ( .A0(n12623), .A1(n12622), .S(n4074), .Z(n12638) );
  CMX2X1 U23076 ( .A0(n12624), .A1(n12638), .S(n3806), .Z(n12647) );
  CMXI2X1 U23077 ( .A0(n12625), .A1(n12647), .S(n3500), .Z(N6145) );
  CMX2X1 U23078 ( .A0(n12627), .A1(n12626), .S(n3807), .Z(n12649) );
  CMXI2X1 U23079 ( .A0(n12628), .A1(n12649), .S(n3501), .Z(N6146) );
  CMX2X1 U23080 ( .A0(n12630), .A1(n12629), .S(n3808), .Z(n12651) );
  CMXI2X1 U23081 ( .A0(n12631), .A1(n12651), .S(n3272), .Z(N6147) );
  CMXI2X1 U23082 ( .A0(n12633), .A1(n12632), .S(n3272), .Z(N5256) );
  CMX2X1 U23083 ( .A0(n12635), .A1(n12634), .S(n3809), .Z(n12653) );
  CMXI2X1 U23084 ( .A0(n12636), .A1(n12653), .S(n3272), .Z(N6148) );
  CMX2X1 U23085 ( .A0(n12638), .A1(n12637), .S(n3797), .Z(n12655) );
  CMXI2X1 U23086 ( .A0(n12639), .A1(n12655), .S(n3272), .Z(N6149) );
  CMXI2X1 U23087 ( .A0(n12641), .A1(n12640), .S(n3272), .Z(N6150) );
  CMXI2X1 U23088 ( .A0(n12643), .A1(n12642), .S(n3272), .Z(N6151) );
  CMXI2X1 U23089 ( .A0(n12645), .A1(n12644), .S(n3272), .Z(N6152) );
  CMXI2X1 U23090 ( .A0(n12647), .A1(n12646), .S(n3272), .Z(N6153) );
  CMXI2X1 U23091 ( .A0(n12649), .A1(n12648), .S(n3272), .Z(N6154) );
  CMXI2X1 U23092 ( .A0(n12651), .A1(n12650), .S(n3272), .Z(N6155) );
  CMXI2X1 U23093 ( .A0(n12653), .A1(n12652), .S(n3272), .Z(N6156) );
  CMXI2X1 U23094 ( .A0(n12655), .A1(n12654), .S(n3273), .Z(N6157) );
  CMXI2X1 U23095 ( .A0(n12657), .A1(n12656), .S(n3273), .Z(N5257) );
  CMXI2X1 U23096 ( .A0(n12659), .A1(n12658), .S(n3273), .Z(N5167) );
  CMXI2X1 U23097 ( .A0(n13400), .A1(n13403), .S(n4202), .Z(n14074) );
  CMXI2X1 U23098 ( .A0(N8277), .A1(N8276), .S(n3879), .Z(n13402) );
  CMXI2X1 U23099 ( .A0(N8278), .A1(N8279), .S(n3889), .Z(n12660) );
  CMXI2X1 U23100 ( .A0(n13402), .A1(n12660), .S(n4202), .Z(n12661) );
  CMXI2X1 U23101 ( .A0(n14074), .A1(n12661), .S(n3778), .Z(n12662) );
  CMX2X1 U23102 ( .A0(N8269), .A1(N8268), .S(n3862), .Z(n12757) );
  CMXI2X1 U23103 ( .A0(N8270), .A1(N8271), .S(n3883), .Z(n13401) );
  CMXI2X1 U23104 ( .A0(n12757), .A1(n4432), .S(n4201), .Z(n14073) );
  CMX2X1 U23105 ( .A0(N8265), .A1(N8264), .S(n3877), .Z(n12759) );
  CMX2X1 U23106 ( .A0(N8267), .A1(N8266), .S(n3863), .Z(n12758) );
  CMXI2X1 U23107 ( .A0(n12759), .A1(n12758), .S(n4201), .Z(n12822) );
  CMX2X1 U23108 ( .A0(n14073), .A1(n12822), .S(n3776), .Z(n15412) );
  CMXI2X1 U23109 ( .A0(n12662), .A1(n15412), .S(n3273), .Z(N8280) );
  CMX2X1 U23110 ( .A0(N7277), .A1(N7276), .S(n3879), .Z(n12663) );
  CMXI2X1 U23111 ( .A0(n12663), .A1(n15690), .S(n4201), .Z(n15697) );
  CMX2X1 U23112 ( .A0(N7275), .A1(N7274), .S(n3871), .Z(n12664) );
  CMXI2X1 U23113 ( .A0(n12665), .A1(n12664), .S(n4201), .Z(n12678) );
  CMX2X1 U23114 ( .A0(n15697), .A1(n12678), .S(n3777), .Z(n15711) );
  CMX2X1 U23115 ( .A0(N7271), .A1(N7270), .S(n3862), .Z(n12666) );
  CMXI2X1 U23116 ( .A0(n12667), .A1(n12666), .S(n4201), .Z(n12677) );
  CMX2X1 U23117 ( .A0(N7267), .A1(N7266), .S(n3863), .Z(n12668) );
  CMXI2X1 U23118 ( .A0(n12669), .A1(n12668), .S(n4201), .Z(n12680) );
  CMX2X1 U23119 ( .A0(n12677), .A1(n12680), .S(n3790), .Z(n12695) );
  CMXI2X1 U23120 ( .A0(n15711), .A1(n12695), .S(n3271), .Z(N9280) );
  CMX2X1 U23121 ( .A0(N7276), .A1(N7275), .S(n3864), .Z(n12670) );
  CMX2X1 U23122 ( .A0(N7278), .A1(N7277), .S(n3865), .Z(n15694) );
  CMXI2X1 U23123 ( .A0(n12670), .A1(n15694), .S(n4201), .Z(n15700) );
  CMX2X1 U23124 ( .A0(N7274), .A1(N7273), .S(n3875), .Z(n12671) );
  CMXI2X1 U23125 ( .A0(n12672), .A1(n12671), .S(n4201), .Z(n12682) );
  CMX2X1 U23126 ( .A0(n15700), .A1(n12682), .S(n3791), .Z(n15713) );
  CMX2X1 U23127 ( .A0(N7268), .A1(N7267), .S(n3876), .Z(n12674) );
  CMXI2X1 U23128 ( .A0(n12674), .A1(n12673), .S(n4201), .Z(n12681) );
  CMX2X1 U23129 ( .A0(N7264), .A1(N7263), .S(n3866), .Z(n12676) );
  CMXI2X1 U23130 ( .A0(n12676), .A1(n12675), .S(n4201), .Z(n12684) );
  CMX2X1 U23131 ( .A0(n12681), .A1(n12684), .S(n3792), .Z(n12698) );
  CMXI2X1 U23132 ( .A0(n15713), .A1(n12698), .S(n3271), .Z(N9281) );
  CMXI2X1 U23133 ( .A0(n12664), .A1(n12663), .S(n4201), .Z(n15705) );
  CMXI2X1 U23134 ( .A0(n12666), .A1(n12665), .S(n4201), .Z(n12686) );
  CMX2X1 U23135 ( .A0(n15705), .A1(n12686), .S(n3793), .Z(n15715) );
  CMXI2X1 U23136 ( .A0(n12668), .A1(n12667), .S(n4201), .Z(n12685) );
  CMX2X1 U23137 ( .A0(N7263), .A1(N7262), .S(n3871), .Z(n12679) );
  CMXI2X1 U23138 ( .A0(n12679), .A1(n12669), .S(n4201), .Z(n12688) );
  CMX2X1 U23139 ( .A0(n12685), .A1(n12688), .S(n3794), .Z(n12701) );
  CMXI2X1 U23140 ( .A0(n15715), .A1(n12701), .S(n3271), .Z(N9282) );
  CMXI2X1 U23141 ( .A0(n12671), .A1(n12670), .S(n4201), .Z(n15708) );
  CMXI2X1 U23142 ( .A0(n12673), .A1(n12672), .S(n4201), .Z(n12690) );
  CMX2X1 U23143 ( .A0(n15708), .A1(n12690), .S(n3795), .Z(n15717) );
  CMXI2X1 U23144 ( .A0(n12675), .A1(n12674), .S(n4200), .Z(n12689) );
  CMXI2X1 U23145 ( .A0(n12683), .A1(n12676), .S(n4200), .Z(n12692) );
  CMX2X1 U23146 ( .A0(n12689), .A1(n12692), .S(n3796), .Z(n12704) );
  CMXI2X1 U23147 ( .A0(n15717), .A1(n12704), .S(n3271), .Z(N9283) );
  CMX2X1 U23148 ( .A0(n12678), .A1(n12677), .S(n3797), .Z(n15719) );
  CMXI2X1 U23149 ( .A0(n12687), .A1(n12679), .S(n4200), .Z(n12694) );
  CMX2X1 U23150 ( .A0(n12680), .A1(n12694), .S(n3805), .Z(n12706) );
  CMXI2X1 U23151 ( .A0(n15719), .A1(n12706), .S(n3271), .Z(N9284) );
  CMX2X1 U23152 ( .A0(n12682), .A1(n12681), .S(n3806), .Z(n15721) );
  CMX2X1 U23153 ( .A0(N7260), .A1(N7259), .S(n3869), .Z(n12691) );
  CMXI2X1 U23154 ( .A0(n12691), .A1(n12683), .S(n4200), .Z(n12697) );
  CMX2X1 U23155 ( .A0(n12684), .A1(n12697), .S(n3790), .Z(n12708) );
  CMXI2X1 U23156 ( .A0(n15721), .A1(n12708), .S(n3271), .Z(N9285) );
  CMX2X1 U23157 ( .A0(n12686), .A1(n12685), .S(n4305), .Z(n15723) );
  CMXI2X1 U23158 ( .A0(n12693), .A1(n12687), .S(n4200), .Z(n12700) );
  CMX2X1 U23159 ( .A0(n12688), .A1(n12700), .S(n3775), .Z(n12710) );
  CMX2X1 U23160 ( .A0(n12690), .A1(n12689), .S(n3776), .Z(n15725) );
  CMX2X1 U23161 ( .A0(N7258), .A1(N7257), .S(n3867), .Z(n12696) );
  CMXI2X1 U23162 ( .A0(n12696), .A1(n12691), .S(n4200), .Z(n12703) );
  CMX2X1 U23163 ( .A0(n12692), .A1(n12703), .S(n3777), .Z(n12712) );
  CMXI2X1 U23164 ( .A0(n12699), .A1(n12693), .S(n4200), .Z(n12705) );
  CMX2X1 U23165 ( .A0(n12694), .A1(n12705), .S(n3807), .Z(n12713) );
  CMXI2X1 U23166 ( .A0(n12695), .A1(n12713), .S(n3271), .Z(N9288) );
  CMXI2X1 U23167 ( .A0(n12702), .A1(n12696), .S(n4200), .Z(n12707) );
  CMX2X1 U23168 ( .A0(n12697), .A1(n12707), .S(n3808), .Z(n12714) );
  CMXI2X1 U23169 ( .A0(n12698), .A1(n12714), .S(n3523), .Z(N9289) );
  CMX2X1 U23170 ( .A0(N8177), .A1(N8176), .S(n3864), .Z(n12721) );
  CMX2X1 U23171 ( .A0(N8179), .A1(N8178), .S(n3865), .Z(n15308) );
  CMXI2X1 U23172 ( .A0(n12721), .A1(n15308), .S(n4200), .Z(n15375) );
  CMX2X1 U23173 ( .A0(N8173), .A1(N8172), .S(n3873), .Z(n12723) );
  CMX2X1 U23174 ( .A0(N8175), .A1(N8174), .S(n3867), .Z(n12722) );
  CMXI2X1 U23175 ( .A0(n12723), .A1(n12722), .S(n4200), .Z(n12736) );
  CMX2X1 U23176 ( .A0(n15375), .A1(n12736), .S(n3790), .Z(n15509) );
  CMX2X1 U23177 ( .A0(N8169), .A1(N8168), .S(n3868), .Z(n12725) );
  CMX2X1 U23178 ( .A0(N8171), .A1(N8170), .S(n3869), .Z(n12724) );
  CMXI2X1 U23179 ( .A0(n12725), .A1(n12724), .S(n4200), .Z(n12735) );
  CMX2X1 U23180 ( .A0(N8165), .A1(N8164), .S(n3873), .Z(n12727) );
  CMX2X1 U23181 ( .A0(N8167), .A1(N8166), .S(n3874), .Z(n12726) );
  CMXI2X1 U23182 ( .A0(n12727), .A1(n12726), .S(n4200), .Z(n12738) );
  CMX2X1 U23183 ( .A0(n12735), .A1(n12738), .S(n3791), .Z(n12753) );
  CMXI2X1 U23184 ( .A0(n15509), .A1(n12753), .S(n3524), .Z(N8380) );
  CMX2X1 U23185 ( .A0(n12700), .A1(n12709), .S(n3809), .Z(n12715) );
  CMXI2X1 U23186 ( .A0(n12701), .A1(n12715), .S(n3520), .Z(N9290) );
  CMX2X1 U23187 ( .A0(n12703), .A1(n12711), .S(n3810), .Z(n12716) );
  CMXI2X1 U23188 ( .A0(n12704), .A1(n12716), .S(n3271), .Z(N9291) );
  CMXI2X1 U23189 ( .A0(n12706), .A1(n12717), .S(n3519), .Z(N9292) );
  CMXI2X1 U23190 ( .A0(n12708), .A1(n12718), .S(n3522), .Z(N9293) );
  CMX2X1 U23191 ( .A0(N8176), .A1(N8175), .S(n3871), .Z(n12728) );
  CMX2X1 U23192 ( .A0(N8178), .A1(N8177), .S(n3866), .Z(n15342) );
  CMXI2X1 U23193 ( .A0(n12728), .A1(n15342), .S(n4200), .Z(n15408) );
  CMX2X1 U23194 ( .A0(N8172), .A1(N8171), .S(n3867), .Z(n12730) );
  CMX2X1 U23195 ( .A0(N8174), .A1(N8173), .S(n3868), .Z(n12729) );
  CMXI2X1 U23196 ( .A0(n12730), .A1(n12729), .S(n4200), .Z(n12740) );
  CMX2X1 U23197 ( .A0(n15408), .A1(n12740), .S(n3797), .Z(n15541) );
  CMX2X1 U23198 ( .A0(N8168), .A1(N8167), .S(n3869), .Z(n12732) );
  CMX2X1 U23199 ( .A0(N8170), .A1(N8169), .S(n3870), .Z(n12731) );
  CMXI2X1 U23200 ( .A0(n12732), .A1(n12731), .S(n4200), .Z(n12739) );
  CMX2X1 U23201 ( .A0(N8164), .A1(N8163), .S(n3879), .Z(n12734) );
  CMX2X1 U23202 ( .A0(N8166), .A1(N8165), .S(n3880), .Z(n12733) );
  CMXI2X1 U23203 ( .A0(n12734), .A1(n12733), .S(n4200), .Z(n12742) );
  CMX2X1 U23204 ( .A0(n12739), .A1(n12742), .S(n3807), .Z(n12756) );
  CMXI2X1 U23205 ( .A0(n15541), .A1(n12756), .S(n3521), .Z(N8381) );
  CMXI2X1 U23206 ( .A0(n12722), .A1(n12721), .S(n4199), .Z(n15443) );
  CMXI2X1 U23207 ( .A0(n12724), .A1(n12723), .S(n4199), .Z(n12744) );
  CMX2X1 U23208 ( .A0(n15443), .A1(n12744), .S(n3808), .Z(n15573) );
  CMX2X1 U23209 ( .A0(N8163), .A1(N8162), .S(n3881), .Z(n12737) );
  CMXI2X1 U23210 ( .A0(n12737), .A1(n12727), .S(n4199), .Z(n12746) );
  CMX2X1 U23211 ( .A0(n12743), .A1(n12746), .S(n3809), .Z(n12762) );
  CMXI2X1 U23212 ( .A0(n15573), .A1(n12762), .S(n3278), .Z(N8382) );
  CMXI2X1 U23213 ( .A0(n12729), .A1(n12728), .S(n4199), .Z(n15476) );
  CMXI2X1 U23214 ( .A0(n12731), .A1(n12730), .S(n4199), .Z(n12748) );
  CMX2X1 U23215 ( .A0(n15476), .A1(n12748), .S(n3810), .Z(n15605) );
  CMX2X1 U23216 ( .A0(N8162), .A1(N8161), .S(n3872), .Z(n12741) );
  CMXI2X1 U23217 ( .A0(n12741), .A1(n12734), .S(n4199), .Z(n12750) );
  CMX2X1 U23218 ( .A0(n12747), .A1(n12750), .S(n3811), .Z(n12765) );
  CMXI2X1 U23219 ( .A0(n15605), .A1(n12765), .S(n3278), .Z(N8383) );
  CMX2X1 U23220 ( .A0(n12736), .A1(n12735), .S(n3812), .Z(n15637) );
  CMX2X1 U23221 ( .A0(N8161), .A1(N8160), .S(n3874), .Z(n12745) );
  CMXI2X1 U23222 ( .A0(n12745), .A1(n12737), .S(n4199), .Z(n12752) );
  CMX2X1 U23223 ( .A0(n12738), .A1(n12752), .S(n4374), .Z(n12768) );
  CMXI2X1 U23224 ( .A0(n15637), .A1(n12768), .S(n3278), .Z(N8384) );
  CMX2X1 U23225 ( .A0(n12740), .A1(n12739), .S(n3771), .Z(n15669) );
  CMX2X1 U23226 ( .A0(N8160), .A1(N8159), .S(n3873), .Z(n12749) );
  CMX2X1 U23227 ( .A0(n12742), .A1(n12755), .S(n3772), .Z(n12771) );
  CMXI2X1 U23228 ( .A0(n15669), .A1(n12771), .S(n3278), .Z(N8385) );
  CMX2X1 U23229 ( .A0(n12744), .A1(n12743), .S(n3773), .Z(n15703) );
  CMX2X1 U23230 ( .A0(N8159), .A1(N8158), .S(n3874), .Z(n12751) );
  CMX2X1 U23231 ( .A0(n12746), .A1(n12761), .S(n3774), .Z(n12774) );
  CMXI2X1 U23232 ( .A0(n15703), .A1(n12774), .S(n3278), .Z(N8386) );
  CMX2X1 U23233 ( .A0(n12748), .A1(n12747), .S(n3775), .Z(n15727) );
  CMX2X1 U23234 ( .A0(N8158), .A1(N8157), .S(n3870), .Z(n12754) );
  CMXI2X1 U23235 ( .A0(n12754), .A1(n12749), .S(n4199), .Z(n12764) );
  CMX2X1 U23236 ( .A0(n12750), .A1(n12764), .S(n3776), .Z(n12777) );
  CMXI2X1 U23237 ( .A0(n15727), .A1(n12777), .S(n3278), .Z(N8387) );
  CMX2X1 U23238 ( .A0(N8157), .A1(N8156), .S(n3876), .Z(n12760) );
  CMX2X1 U23239 ( .A0(n12752), .A1(n12767), .S(n3777), .Z(n12780) );
  CMXI2X1 U23240 ( .A0(n12753), .A1(n12780), .S(n3278), .Z(N8388) );
  CMX2X1 U23241 ( .A0(N8156), .A1(N8155), .S(n3877), .Z(n12763) );
  CMXI2X1 U23242 ( .A0(n12763), .A1(n12754), .S(n4199), .Z(n12770) );
  CMX2X1 U23243 ( .A0(n12755), .A1(n12770), .S(n3790), .Z(n12783) );
  CMXI2X1 U23244 ( .A0(n12756), .A1(n12783), .S(n3278), .Z(N8389) );
  CMXI2X1 U23245 ( .A0(n12758), .A1(n12757), .S(n4199), .Z(n14741) );
  CMX2X1 U23246 ( .A0(N8263), .A1(N8262), .S(n3878), .Z(n12820) );
  CMXI2X1 U23247 ( .A0(n12820), .A1(n12759), .S(n4199), .Z(n12894) );
  CMX2X1 U23248 ( .A0(n14741), .A1(n12894), .S(n3791), .Z(n13405) );
  CMX2X1 U23249 ( .A0(N8259), .A1(N8258), .S(n3862), .Z(n12823) );
  CMX2X1 U23250 ( .A0(N8261), .A1(N8260), .S(n3875), .Z(n12821) );
  CMXI2X1 U23251 ( .A0(n12823), .A1(n12821), .S(n4198), .Z(n12893) );
  CMX2X1 U23252 ( .A0(N8255), .A1(N8254), .S(n3876), .Z(n12825) );
  CMX2X1 U23253 ( .A0(N8257), .A1(N8256), .S(n3870), .Z(n12824) );
  CMXI2X1 U23254 ( .A0(n12825), .A1(n12824), .S(n4198), .Z(n12896) );
  CMX2X1 U23255 ( .A0(n12893), .A1(n12896), .S(n3791), .Z(n13031) );
  CMXI2X1 U23256 ( .A0(n13405), .A1(n13031), .S(n3278), .Z(N8290) );
  CMX2X1 U23257 ( .A0(N8155), .A1(N8154), .S(n3875), .Z(n12766) );
  CMXI2X1 U23258 ( .A0(n12766), .A1(n12760), .S(n4198), .Z(n12773) );
  CMX2X1 U23259 ( .A0(n12761), .A1(n12773), .S(n3810), .Z(n12786) );
  CMX2X1 U23260 ( .A0(N8154), .A1(N8153), .S(n3871), .Z(n12769) );
  CMX2X1 U23261 ( .A0(n12764), .A1(n12776), .S(n3811), .Z(n12789) );
  CMXI2X1 U23262 ( .A0(n12765), .A1(n12789), .S(n3277), .Z(N8391) );
  CMX2X1 U23263 ( .A0(N8153), .A1(N8152), .S(n3880), .Z(n12772) );
  CMXI2X1 U23264 ( .A0(n12772), .A1(n12766), .S(n4198), .Z(n12779) );
  CMX2X1 U23265 ( .A0(n3711), .A1(n12779), .S(n3812), .Z(n12792) );
  CMXI2X1 U23266 ( .A0(n12768), .A1(n12792), .S(n3277), .Z(N8392) );
  CMX2X1 U23267 ( .A0(N8152), .A1(N8151), .S(n3879), .Z(n12775) );
  CMX2X1 U23268 ( .A0(n12770), .A1(n12782), .S(n4306), .Z(n12795) );
  CMXI2X1 U23269 ( .A0(n12771), .A1(n12795), .S(n3273), .Z(N8393) );
  CMX2X1 U23270 ( .A0(N8151), .A1(N8150), .S(n3869), .Z(n12778) );
  CMXI2X1 U23271 ( .A0(n12778), .A1(n12772), .S(n4198), .Z(n12785) );
  CMX2X1 U23272 ( .A0(n12773), .A1(n12785), .S(n3771), .Z(n12798) );
  CMX2X1 U23273 ( .A0(N8150), .A1(N8149), .S(n3868), .Z(n12781) );
  CMXI2X1 U23274 ( .A0(n12781), .A1(n12775), .S(n4198), .Z(n12788) );
  CMX2X1 U23275 ( .A0(n12776), .A1(n12788), .S(n3795), .Z(n12801) );
  CMXI2X1 U23276 ( .A0(n12777), .A1(n12801), .S(n3439), .Z(N8395) );
  CMX2X1 U23277 ( .A0(N8149), .A1(N8148), .S(n3876), .Z(n12784) );
  CMXI2X1 U23278 ( .A0(n12784), .A1(n12778), .S(n4198), .Z(n12791) );
  CMX2X1 U23279 ( .A0(n12779), .A1(n12791), .S(n3772), .Z(n12804) );
  CMX2X1 U23280 ( .A0(N8148), .A1(N8147), .S(n3877), .Z(n12787) );
  CMXI2X1 U23281 ( .A0(n12787), .A1(n12781), .S(n4198), .Z(n12794) );
  CMX2X1 U23282 ( .A0(n12782), .A1(n12794), .S(n3806), .Z(n12807) );
  CMX2X1 U23283 ( .A0(N8147), .A1(N8146), .S(n3869), .Z(n12790) );
  CMXI2X1 U23284 ( .A0(n12790), .A1(n12784), .S(n4198), .Z(n12797) );
  CMX2X1 U23285 ( .A0(n12785), .A1(n12797), .S(n3807), .Z(n12810) );
  CMXI2X1 U23286 ( .A0(n12786), .A1(n12810), .S(n3271), .Z(N8398) );
  CMX2X1 U23287 ( .A0(N8146), .A1(N8145), .S(n3870), .Z(n12793) );
  CMXI2X1 U23288 ( .A0(n12793), .A1(n12787), .S(n4198), .Z(n12800) );
  CMX2X1 U23289 ( .A0(n12788), .A1(n12800), .S(n3808), .Z(n12813) );
  CMXI2X1 U23290 ( .A0(n12789), .A1(n12813), .S(n3280), .Z(N8399) );
  CMX2X1 U23291 ( .A0(N8266), .A1(N8265), .S(n3866), .Z(n12856) );
  CMX2X1 U23292 ( .A0(N8268), .A1(N8267), .S(n3865), .Z(n13067) );
  CMXI2X1 U23293 ( .A0(n12856), .A1(n13067), .S(n4198), .Z(n15075) );
  CMX2X1 U23294 ( .A0(N8262), .A1(N8261), .S(n3877), .Z(n12858) );
  CMX2X1 U23295 ( .A0(N8264), .A1(N8263), .S(n3878), .Z(n12857) );
  CMXI2X1 U23296 ( .A0(n12858), .A1(n12857), .S(n4198), .Z(n12928) );
  CMX2X1 U23297 ( .A0(n15075), .A1(n12928), .S(n3809), .Z(n13742) );
  CMX2X1 U23298 ( .A0(N8258), .A1(N8257), .S(n3879), .Z(n12860) );
  CMX2X1 U23299 ( .A0(N8260), .A1(N8259), .S(n3880), .Z(n12859) );
  CMXI2X1 U23300 ( .A0(n12860), .A1(n12859), .S(n4198), .Z(n12927) );
  CMX2X1 U23301 ( .A0(N8254), .A1(N8253), .S(n3875), .Z(n12862) );
  CMX2X1 U23302 ( .A0(N8256), .A1(N8255), .S(n3876), .Z(n12861) );
  CMXI2X1 U23303 ( .A0(n12862), .A1(n12861), .S(n4198), .Z(n12930) );
  CMX2X1 U23304 ( .A0(n12927), .A1(n12930), .S(n3793), .Z(n13064) );
  CMXI2X1 U23305 ( .A0(n13742), .A1(n13064), .S(n3280), .Z(N8291) );
  CMX2X1 U23306 ( .A0(N8145), .A1(N8144), .S(n3877), .Z(n12796) );
  CMXI2X1 U23307 ( .A0(n12796), .A1(n12790), .S(n4197), .Z(n12803) );
  CMX2X1 U23308 ( .A0(n12791), .A1(n12803), .S(n3794), .Z(n12816) );
  CMXI2X1 U23309 ( .A0(n12792), .A1(n12816), .S(n3280), .Z(N8400) );
  CMX2X1 U23310 ( .A0(N8144), .A1(N8143), .S(n3878), .Z(n12799) );
  CMXI2X1 U23311 ( .A0(n12799), .A1(n12793), .S(n4197), .Z(n12806) );
  CMX2X1 U23312 ( .A0(n12794), .A1(n12806), .S(n3795), .Z(n12819) );
  CMXI2X1 U23313 ( .A0(n12795), .A1(n12819), .S(n3280), .Z(N8401) );
  CMX2X1 U23314 ( .A0(N8143), .A1(N8142), .S(n3875), .Z(n12802) );
  CMXI2X1 U23315 ( .A0(n12802), .A1(n12796), .S(n4197), .Z(n12809) );
  CMX2X1 U23316 ( .A0(n12797), .A1(n12809), .S(n3796), .Z(n12828) );
  CMXI2X1 U23317 ( .A0(n12798), .A1(n12828), .S(n3280), .Z(N8402) );
  CMX2X1 U23318 ( .A0(N8142), .A1(N8141), .S(n3871), .Z(n12805) );
  CMXI2X1 U23319 ( .A0(n12805), .A1(n12799), .S(n4197), .Z(n12812) );
  CMX2X1 U23320 ( .A0(n12800), .A1(n12812), .S(n3797), .Z(n12831) );
  CMXI2X1 U23321 ( .A0(n12801), .A1(n12831), .S(n3279), .Z(N8403) );
  CMX2X1 U23322 ( .A0(N8141), .A1(N8140), .S(n3872), .Z(n12808) );
  CMXI2X1 U23323 ( .A0(n12808), .A1(n12802), .S(n4197), .Z(n12815) );
  CMX2X1 U23324 ( .A0(n12803), .A1(n12815), .S(n3805), .Z(n12834) );
  CMXI2X1 U23325 ( .A0(n12804), .A1(n12834), .S(n3279), .Z(N8404) );
  CMX2X1 U23326 ( .A0(N8140), .A1(N8139), .S(n3873), .Z(n12811) );
  CMXI2X1 U23327 ( .A0(n12811), .A1(n12805), .S(n4197), .Z(n12818) );
  CMX2X1 U23328 ( .A0(n12806), .A1(n12818), .S(n3806), .Z(n12837) );
  CMXI2X1 U23329 ( .A0(n12807), .A1(n12837), .S(n3279), .Z(N8405) );
  CMX2X1 U23330 ( .A0(N8139), .A1(N8138), .S(n3874), .Z(n12814) );
  CMXI2X1 U23331 ( .A0(n12814), .A1(n12808), .S(n4197), .Z(n12827) );
  CMX2X1 U23332 ( .A0(n12809), .A1(n12827), .S(n3807), .Z(n12840) );
  CMXI2X1 U23333 ( .A0(n12810), .A1(n12840), .S(n3279), .Z(N8406) );
  CMX2X1 U23334 ( .A0(N8138), .A1(N8137), .S(n3875), .Z(n12817) );
  CMXI2X1 U23335 ( .A0(n12817), .A1(n12811), .S(n4197), .Z(n12830) );
  CMX2X1 U23336 ( .A0(n12812), .A1(n12830), .S(n3808), .Z(n12843) );
  CMXI2X1 U23337 ( .A0(n12813), .A1(n12843), .S(n3279), .Z(N8407) );
  CMX2X1 U23338 ( .A0(N8137), .A1(N8136), .S(n3876), .Z(n12826) );
  CMXI2X1 U23339 ( .A0(n12826), .A1(n12814), .S(n4197), .Z(n12833) );
  CMX2X1 U23340 ( .A0(n12815), .A1(n12833), .S(n3775), .Z(n12846) );
  CMXI2X1 U23341 ( .A0(n12816), .A1(n12846), .S(n3279), .Z(N8408) );
  CMX2X1 U23342 ( .A0(N8136), .A1(N8135), .S(n3877), .Z(n12829) );
  CMXI2X1 U23343 ( .A0(n12829), .A1(n12817), .S(n4197), .Z(n12836) );
  CMX2X1 U23344 ( .A0(n12818), .A1(n12836), .S(n3772), .Z(n12849) );
  CMXI2X1 U23345 ( .A0(n12819), .A1(n12849), .S(n3279), .Z(N8409) );
  CMXI2X1 U23346 ( .A0(n12821), .A1(n12820), .S(n4197), .Z(n12962) );
  CMX2X1 U23347 ( .A0(n12822), .A1(n12962), .S(n3773), .Z(n14075) );
  CMXI2X1 U23348 ( .A0(n12824), .A1(n12823), .S(n4197), .Z(n12961) );
  CMX2X1 U23349 ( .A0(N8253), .A1(N8252), .S(n3878), .Z(n12895) );
  CMXI2X1 U23350 ( .A0(n12895), .A1(n12825), .S(n4197), .Z(n12964) );
  CMX2X1 U23351 ( .A0(n12961), .A1(n12964), .S(n3774), .Z(n13102) );
  CMXI2X1 U23352 ( .A0(n14075), .A1(n13102), .S(n3279), .Z(N8292) );
  CMX2X1 U23353 ( .A0(N8135), .A1(N8134), .S(n3879), .Z(n12832) );
  CMXI2X1 U23354 ( .A0(n12832), .A1(n12826), .S(n4197), .Z(n12839) );
  CMX2X1 U23355 ( .A0(n12827), .A1(n12839), .S(n3775), .Z(n12852) );
  CMXI2X1 U23356 ( .A0(n12828), .A1(n12852), .S(n3279), .Z(N8410) );
  CMX2X1 U23357 ( .A0(N8134), .A1(N8133), .S(n3878), .Z(n12835) );
  CMXI2X1 U23358 ( .A0(n12835), .A1(n12829), .S(n4197), .Z(n12842) );
  CMX2X1 U23359 ( .A0(n12830), .A1(n12842), .S(n3808), .Z(n12855) );
  CMXI2X1 U23360 ( .A0(n12831), .A1(n12855), .S(n3279), .Z(N8411) );
  CMX2X1 U23361 ( .A0(N8133), .A1(N8132), .S(n3879), .Z(n12838) );
  CMXI2X1 U23362 ( .A0(n12838), .A1(n12832), .S(n4197), .Z(n12845) );
  CMX2X1 U23363 ( .A0(n12833), .A1(n12845), .S(n3792), .Z(n12865) );
  CMXI2X1 U23364 ( .A0(n12834), .A1(n12865), .S(n3279), .Z(N8412) );
  CMX2X1 U23365 ( .A0(N8132), .A1(N8131), .S(n3881), .Z(n12841) );
  CMXI2X1 U23366 ( .A0(n12841), .A1(n12835), .S(n4196), .Z(n12848) );
  CMX2X1 U23367 ( .A0(n12836), .A1(n12848), .S(n3793), .Z(n12868) );
  CMXI2X1 U23368 ( .A0(n12837), .A1(n12868), .S(n3278), .Z(N8413) );
  CMX2X1 U23369 ( .A0(N8131), .A1(N8130), .S(n3862), .Z(n12844) );
  CMXI2X1 U23370 ( .A0(n12844), .A1(n12838), .S(n4196), .Z(n12851) );
  CMX2X1 U23371 ( .A0(n12839), .A1(n12851), .S(n3794), .Z(n12871) );
  CMXI2X1 U23372 ( .A0(n12840), .A1(n12871), .S(n3278), .Z(N8414) );
  CMX2X1 U23373 ( .A0(N8130), .A1(N8129), .S(n3863), .Z(n12847) );
  CMXI2X1 U23374 ( .A0(n12847), .A1(n12841), .S(n4196), .Z(n12854) );
  CMX2X1 U23375 ( .A0(n12842), .A1(n12854), .S(n3795), .Z(n12874) );
  CMXI2X1 U23376 ( .A0(n12843), .A1(n12874), .S(n3292), .Z(N8415) );
  CMX2X1 U23377 ( .A0(N8129), .A1(N8128), .S(n3864), .Z(n12850) );
  CMXI2X1 U23378 ( .A0(n12850), .A1(n12844), .S(n4196), .Z(n12864) );
  CMX2X1 U23379 ( .A0(n12845), .A1(n12864), .S(n3796), .Z(n12877) );
  CMXI2X1 U23380 ( .A0(n12846), .A1(n12877), .S(n3492), .Z(N8416) );
  CMX2X1 U23381 ( .A0(N8128), .A1(N8127), .S(n3879), .Z(n12853) );
  CMXI2X1 U23382 ( .A0(n12853), .A1(n12847), .S(n4196), .Z(n12867) );
  CMX2X1 U23383 ( .A0(n12848), .A1(n12867), .S(n3797), .Z(n12880) );
  CMXI2X1 U23384 ( .A0(n12849), .A1(n12880), .S(n3491), .Z(N8417) );
  CMX2X1 U23385 ( .A0(N8127), .A1(N8126), .S(n3880), .Z(n12863) );
  CMXI2X1 U23386 ( .A0(n12863), .A1(n12850), .S(n4196), .Z(n12870) );
  CMX2X1 U23387 ( .A0(n12851), .A1(n12870), .S(n3805), .Z(n12883) );
  CMXI2X1 U23388 ( .A0(n12852), .A1(n12883), .S(n3490), .Z(N8418) );
  CMX2X1 U23389 ( .A0(N8126), .A1(N8125), .S(n3881), .Z(n12866) );
  CMXI2X1 U23390 ( .A0(n12866), .A1(n12853), .S(n4196), .Z(n12873) );
  CMX2X1 U23391 ( .A0(n12854), .A1(n12873), .S(n3806), .Z(n12886) );
  CMXI2X1 U23392 ( .A0(n12855), .A1(n12886), .S(n3489), .Z(N8419) );
  CMXI2X1 U23393 ( .A0(n12857), .A1(n12856), .S(n4196), .Z(n13068) );
  CMXI2X1 U23394 ( .A0(n12859), .A1(n12858), .S(n4196), .Z(n12996) );
  CMX2X1 U23395 ( .A0(n13068), .A1(n12996), .S(n3807), .Z(n14409) );
  CMXI2X1 U23396 ( .A0(n12861), .A1(n12860), .S(n4196), .Z(n12995) );
  CMX2X1 U23397 ( .A0(N8252), .A1(N8251), .S(n3862), .Z(n12929) );
  CMXI2X1 U23398 ( .A0(n12929), .A1(n12862), .S(n4196), .Z(n12998) );
  CMX2X1 U23399 ( .A0(n12995), .A1(n12998), .S(n3808), .Z(n13135) );
  CMXI2X1 U23400 ( .A0(n14409), .A1(n13135), .S(n3488), .Z(N8293) );
  CMX2X1 U23401 ( .A0(N8125), .A1(N8124), .S(n3876), .Z(n12869) );
  CMXI2X1 U23402 ( .A0(n12869), .A1(n12863), .S(n4196), .Z(n12876) );
  CMX2X1 U23403 ( .A0(n12864), .A1(n12876), .S(n3809), .Z(n12889) );
  CMXI2X1 U23404 ( .A0(n12865), .A1(n12889), .S(n3487), .Z(N8420) );
  CMX2X1 U23405 ( .A0(N8124), .A1(N8123), .S(n3880), .Z(n12872) );
  CMXI2X1 U23406 ( .A0(n12872), .A1(n12866), .S(n4196), .Z(n12879) );
  CMX2X1 U23407 ( .A0(n12867), .A1(n12879), .S(n3810), .Z(n12892) );
  CMXI2X1 U23408 ( .A0(n12868), .A1(n12892), .S(n3288), .Z(N8421) );
  CMX2X1 U23409 ( .A0(N8123), .A1(N8122), .S(n3881), .Z(n12875) );
  CMXI2X1 U23410 ( .A0(n12875), .A1(n12869), .S(n4196), .Z(n12882) );
  CMX2X1 U23411 ( .A0(n12870), .A1(n12882), .S(n3811), .Z(n12899) );
  CMXI2X1 U23412 ( .A0(n12871), .A1(n12899), .S(n3288), .Z(N8422) );
  CMX2X1 U23413 ( .A0(N8122), .A1(N8121), .S(n3862), .Z(n12878) );
  CMXI2X1 U23414 ( .A0(n12878), .A1(n12872), .S(n4196), .Z(n12885) );
  CMX2X1 U23415 ( .A0(n12873), .A1(n12885), .S(n3812), .Z(n12902) );
  CMXI2X1 U23416 ( .A0(n12874), .A1(n12902), .S(n3288), .Z(N8423) );
  CMX2X1 U23417 ( .A0(N8121), .A1(N8120), .S(n3863), .Z(n12881) );
  CMXI2X1 U23418 ( .A0(n12881), .A1(n12875), .S(n4196), .Z(n12888) );
  CMX2X1 U23419 ( .A0(n12876), .A1(n12888), .S(n4370), .Z(n12905) );
  CMXI2X1 U23420 ( .A0(n12877), .A1(n12905), .S(n3288), .Z(N8424) );
  CMX2X1 U23421 ( .A0(N8120), .A1(N8119), .S(n3864), .Z(n12884) );
  CMXI2X1 U23422 ( .A0(n12884), .A1(n12878), .S(n4195), .Z(n12891) );
  CMX2X1 U23423 ( .A0(n12879), .A1(n12891), .S(n3771), .Z(n12908) );
  CMXI2X1 U23424 ( .A0(n12880), .A1(n12908), .S(n3288), .Z(N8425) );
  CMX2X1 U23425 ( .A0(N8119), .A1(N8118), .S(n3865), .Z(n12887) );
  CMXI2X1 U23426 ( .A0(n12887), .A1(n12881), .S(n4195), .Z(n12898) );
  CMX2X1 U23427 ( .A0(n12882), .A1(n12898), .S(n3795), .Z(n12911) );
  CMXI2X1 U23428 ( .A0(n12883), .A1(n12911), .S(n3288), .Z(N8426) );
  CMX2X1 U23429 ( .A0(N8118), .A1(N8117), .S(n3866), .Z(n12890) );
  CMXI2X1 U23430 ( .A0(n12890), .A1(n12884), .S(n4195), .Z(n12901) );
  CMX2X1 U23431 ( .A0(n12885), .A1(n12901), .S(n3775), .Z(n12914) );
  CMXI2X1 U23432 ( .A0(n12886), .A1(n12914), .S(n3288), .Z(N8427) );
  CMX2X1 U23433 ( .A0(N8117), .A1(N8116), .S(n3880), .Z(n12897) );
  CMXI2X1 U23434 ( .A0(n12897), .A1(n12887), .S(n4195), .Z(n12904) );
  CMX2X1 U23435 ( .A0(n12888), .A1(n12904), .S(n3776), .Z(n12917) );
  CMXI2X1 U23436 ( .A0(n12889), .A1(n12917), .S(n3287), .Z(N8428) );
  CMX2X1 U23437 ( .A0(N8116), .A1(N8115), .S(n3881), .Z(n12900) );
  CMXI2X1 U23438 ( .A0(n12900), .A1(n12890), .S(n4195), .Z(n12907) );
  CMX2X1 U23439 ( .A0(n12891), .A1(n12907), .S(n3777), .Z(n12920) );
  CMXI2X1 U23440 ( .A0(n12892), .A1(n12920), .S(n3287), .Z(N8429) );
  CMX2X1 U23441 ( .A0(n12894), .A1(n12893), .S(n3790), .Z(n14743) );
  CMX2X1 U23442 ( .A0(N8251), .A1(N8250), .S(n3867), .Z(n12963) );
  CMXI2X1 U23443 ( .A0(n12963), .A1(n12895), .S(n4195), .Z(n13030) );
  CMX2X1 U23444 ( .A0(n12896), .A1(n13030), .S(n3791), .Z(n13168) );
  CMXI2X1 U23445 ( .A0(n14743), .A1(n13168), .S(n3287), .Z(N8294) );
  CMX2X1 U23446 ( .A0(N8115), .A1(N8114), .S(n3868), .Z(n12903) );
  CMXI2X1 U23447 ( .A0(n12903), .A1(n12897), .S(n4195), .Z(n12910) );
  CMX2X1 U23448 ( .A0(n12898), .A1(n12910), .S(n3792), .Z(n12923) );
  CMXI2X1 U23449 ( .A0(n12899), .A1(n12923), .S(n3287), .Z(N8430) );
  CMX2X1 U23450 ( .A0(N8114), .A1(N8113), .S(n3865), .Z(n12906) );
  CMXI2X1 U23451 ( .A0(n12906), .A1(n12900), .S(n4195), .Z(n12913) );
  CMX2X1 U23452 ( .A0(n12901), .A1(n12913), .S(n3809), .Z(n12926) );
  CMXI2X1 U23453 ( .A0(n12902), .A1(n12926), .S(n3287), .Z(N8431) );
  CMX2X1 U23454 ( .A0(N8113), .A1(N8112), .S(n3866), .Z(n12909) );
  CMXI2X1 U23455 ( .A0(n12909), .A1(n12903), .S(n4195), .Z(n12916) );
  CMX2X1 U23456 ( .A0(n12904), .A1(n12916), .S(n3772), .Z(n12933) );
  CMXI2X1 U23457 ( .A0(n12905), .A1(n12933), .S(n3287), .Z(N8432) );
  CMX2X1 U23458 ( .A0(N8112), .A1(N8111), .S(n3867), .Z(n12912) );
  CMXI2X1 U23459 ( .A0(n12912), .A1(n12906), .S(n4195), .Z(n12919) );
  CMX2X1 U23460 ( .A0(n12907), .A1(n12919), .S(n3773), .Z(n12936) );
  CMXI2X1 U23461 ( .A0(n12908), .A1(n12936), .S(n3287), .Z(N8433) );
  CMX2X1 U23462 ( .A0(N8111), .A1(N8110), .S(n3868), .Z(n12915) );
  CMXI2X1 U23463 ( .A0(n12915), .A1(n12909), .S(n4195), .Z(n12922) );
  CMX2X1 U23464 ( .A0(n12910), .A1(n12922), .S(n3774), .Z(n12939) );
  CMXI2X1 U23465 ( .A0(n12911), .A1(n12939), .S(n3287), .Z(N8434) );
  CMX2X1 U23466 ( .A0(N8110), .A1(N8109), .S(n3863), .Z(n12918) );
  CMXI2X1 U23467 ( .A0(n12918), .A1(n12912), .S(n4195), .Z(n12925) );
  CMX2X1 U23468 ( .A0(n12913), .A1(n12925), .S(n3775), .Z(n12942) );
  CMXI2X1 U23469 ( .A0(n12914), .A1(n12942), .S(n3287), .Z(N8435) );
  CMX2X1 U23470 ( .A0(N8109), .A1(N8108), .S(n3864), .Z(n12921) );
  CMXI2X1 U23471 ( .A0(n12921), .A1(n12915), .S(n4195), .Z(n12932) );
  CMX2X1 U23472 ( .A0(n12916), .A1(n12932), .S(n3776), .Z(n12945) );
  CMXI2X1 U23473 ( .A0(n12917), .A1(n12945), .S(n3287), .Z(N8436) );
  CMX2X1 U23474 ( .A0(N8108), .A1(N8107), .S(n3865), .Z(n12924) );
  CMXI2X1 U23475 ( .A0(n12924), .A1(n12918), .S(n4195), .Z(n12935) );
  CMX2X1 U23476 ( .A0(n12919), .A1(n12935), .S(n3777), .Z(n12948) );
  CMXI2X1 U23477 ( .A0(n12920), .A1(n12948), .S(n3287), .Z(N8437) );
  CMX2X1 U23478 ( .A0(N8107), .A1(N8106), .S(n3864), .Z(n12931) );
  CMXI2X1 U23479 ( .A0(n12931), .A1(n12921), .S(n4195), .Z(n12938) );
  CMX2X1 U23480 ( .A0(n12922), .A1(n12938), .S(n3790), .Z(n12951) );
  CMXI2X1 U23481 ( .A0(n12923), .A1(n12951), .S(n3290), .Z(N8438) );
  CMX2X1 U23482 ( .A0(N8106), .A1(N8105), .S(n3865), .Z(n12934) );
  CMXI2X1 U23483 ( .A0(n12934), .A1(n12924), .S(n4195), .Z(n12941) );
  CMX2X1 U23484 ( .A0(n12925), .A1(n12941), .S(n3791), .Z(n12954) );
  CMXI2X1 U23485 ( .A0(n12926), .A1(n12954), .S(n3290), .Z(N8439) );
  CMX2X1 U23486 ( .A0(n12928), .A1(n12927), .S(n3792), .Z(n15077) );
  CMX2X1 U23487 ( .A0(N8250), .A1(N8249), .S(n3866), .Z(n12997) );
  CMXI2X1 U23488 ( .A0(n12997), .A1(n12929), .S(n4194), .Z(n13063) );
  CMX2X1 U23489 ( .A0(n12930), .A1(n13063), .S(n3793), .Z(n13201) );
  CMXI2X1 U23490 ( .A0(n15077), .A1(n13201), .S(n3290), .Z(N8295) );
  CMX2X1 U23491 ( .A0(N8105), .A1(N8104), .S(n3867), .Z(n12937) );
  CMXI2X1 U23492 ( .A0(n12937), .A1(n12931), .S(n4194), .Z(n12944) );
  CMX2X1 U23493 ( .A0(n12932), .A1(n12944), .S(n3794), .Z(n12957) );
  CMXI2X1 U23494 ( .A0(n12933), .A1(n12957), .S(n3289), .Z(N8440) );
  CMX2X1 U23495 ( .A0(N8104), .A1(N8103), .S(n3868), .Z(n12940) );
  CMXI2X1 U23496 ( .A0(n12940), .A1(n12934), .S(n4194), .Z(n12947) );
  CMX2X1 U23497 ( .A0(n12935), .A1(n12947), .S(n3795), .Z(n12960) );
  CMXI2X1 U23498 ( .A0(n12936), .A1(n12960), .S(n3289), .Z(N8441) );
  CMX2X1 U23499 ( .A0(N8103), .A1(N8102), .S(n3875), .Z(n12943) );
  CMXI2X1 U23500 ( .A0(n12943), .A1(n12937), .S(n4194), .Z(n12950) );
  CMX2X1 U23501 ( .A0(n12938), .A1(n12950), .S(n3796), .Z(n12967) );
  CMXI2X1 U23502 ( .A0(n12939), .A1(n12967), .S(n3289), .Z(N8442) );
  CMX2X1 U23503 ( .A0(N8102), .A1(N8101), .S(n3876), .Z(n12946) );
  CMXI2X1 U23504 ( .A0(n12946), .A1(n12940), .S(n4194), .Z(n12953) );
  CMX2X1 U23505 ( .A0(n12941), .A1(n12953), .S(n3797), .Z(n12970) );
  CMXI2X1 U23506 ( .A0(n12942), .A1(n12970), .S(n3289), .Z(N8443) );
  CMX2X1 U23507 ( .A0(N8101), .A1(N8100), .S(n3869), .Z(n12949) );
  CMXI2X1 U23508 ( .A0(n12949), .A1(n12943), .S(n4194), .Z(n12956) );
  CMX2X1 U23509 ( .A0(n12944), .A1(n12956), .S(n3805), .Z(n12973) );
  CMXI2X1 U23510 ( .A0(n12945), .A1(n12973), .S(n3289), .Z(N8444) );
  CMX2X1 U23511 ( .A0(N8100), .A1(N8099), .S(n3870), .Z(n12952) );
  CMXI2X1 U23512 ( .A0(n12952), .A1(n12946), .S(n4194), .Z(n12959) );
  CMX2X1 U23513 ( .A0(n12947), .A1(n12959), .S(n3806), .Z(n12976) );
  CMXI2X1 U23514 ( .A0(n12948), .A1(n12976), .S(n3289), .Z(N8445) );
  CMX2X1 U23515 ( .A0(N8099), .A1(N8098), .S(n3881), .Z(n12955) );
  CMXI2X1 U23516 ( .A0(n12955), .A1(n12949), .S(n4194), .Z(n12966) );
  CMX2X1 U23517 ( .A0(n12950), .A1(n12966), .S(n3796), .Z(n12979) );
  CMXI2X1 U23518 ( .A0(n12951), .A1(n12979), .S(n3289), .Z(N8446) );
  CMX2X1 U23519 ( .A0(N8098), .A1(N8097), .S(n3862), .Z(n12958) );
  CMXI2X1 U23520 ( .A0(n12958), .A1(n12952), .S(n4194), .Z(n12969) );
  CMX2X1 U23521 ( .A0(n12953), .A1(n12969), .S(n3776), .Z(n12982) );
  CMXI2X1 U23522 ( .A0(n12954), .A1(n12982), .S(n3289), .Z(N8447) );
  CMX2X1 U23523 ( .A0(N8097), .A1(N8096), .S(n3863), .Z(n12965) );
  CMXI2X1 U23524 ( .A0(n12965), .A1(n12955), .S(n4194), .Z(n12972) );
  CMX2X1 U23525 ( .A0(n12956), .A1(n12972), .S(n3793), .Z(n12985) );
  CMXI2X1 U23526 ( .A0(n12957), .A1(n12985), .S(n3289), .Z(N8448) );
  CMX2X1 U23527 ( .A0(N8096), .A1(N8095), .S(n3864), .Z(n12968) );
  CMXI2X1 U23528 ( .A0(n12968), .A1(n12958), .S(n4194), .Z(n12975) );
  CMX2X1 U23529 ( .A0(n12959), .A1(n12975), .S(n3794), .Z(n12988) );
  CMXI2X1 U23530 ( .A0(n12960), .A1(n12988), .S(n3289), .Z(N8449) );
  CMX2X1 U23531 ( .A0(n12962), .A1(n12961), .S(n3795), .Z(n15411) );
  CMX2X1 U23532 ( .A0(N8249), .A1(N8248), .S(n3874), .Z(n13029) );
  CMXI2X1 U23533 ( .A0(n13029), .A1(n12963), .S(n4194), .Z(n13101) );
  CMX2X1 U23534 ( .A0(n12964), .A1(n13101), .S(n3796), .Z(n13234) );
  CMXI2X1 U23535 ( .A0(n15411), .A1(n13234), .S(n3289), .Z(N8296) );
  CMX2X1 U23536 ( .A0(N8095), .A1(N8094), .S(n3875), .Z(n12971) );
  CMXI2X1 U23537 ( .A0(n12971), .A1(n12965), .S(n4194), .Z(n12978) );
  CMX2X1 U23538 ( .A0(n12966), .A1(n12978), .S(n3797), .Z(n12991) );
  CMXI2X1 U23539 ( .A0(n12967), .A1(n12991), .S(n3288), .Z(N8450) );
  CMX2X1 U23540 ( .A0(N8094), .A1(N8093), .S(n3876), .Z(n12974) );
  CMXI2X1 U23541 ( .A0(n12974), .A1(n12968), .S(n4194), .Z(n12981) );
  CMX2X1 U23542 ( .A0(n12969), .A1(n12981), .S(n3810), .Z(n12994) );
  CMXI2X1 U23543 ( .A0(n12970), .A1(n12994), .S(n3288), .Z(N8451) );
  CMX2X1 U23544 ( .A0(N8093), .A1(N8092), .S(n3877), .Z(n12977) );
  CMXI2X1 U23545 ( .A0(n12977), .A1(n12971), .S(n4194), .Z(n12984) );
  CMX2X1 U23546 ( .A0(n12972), .A1(n12984), .S(n3807), .Z(n13001) );
  CMXI2X1 U23547 ( .A0(n12973), .A1(n13001), .S(n3288), .Z(N8452) );
  CMX2X1 U23548 ( .A0(N8092), .A1(N8091), .S(n3869), .Z(n12980) );
  CMXI2X1 U23549 ( .A0(n12980), .A1(n12974), .S(n4194), .Z(n12987) );
  CMX2X1 U23550 ( .A0(n12975), .A1(n12987), .S(n3808), .Z(n13004) );
  CMXI2X1 U23551 ( .A0(n12976), .A1(n13004), .S(n3288), .Z(N8453) );
  CMX2X1 U23552 ( .A0(N8091), .A1(N8090), .S(n3871), .Z(n12983) );
  CMXI2X1 U23553 ( .A0(n12983), .A1(n12977), .S(n4193), .Z(n12990) );
  CMX2X1 U23554 ( .A0(n12978), .A1(n12990), .S(n3809), .Z(n13007) );
  CMXI2X1 U23555 ( .A0(n12979), .A1(n13007), .S(n3470), .Z(N8454) );
  CMX2X1 U23556 ( .A0(N8090), .A1(N8089), .S(n3872), .Z(n12986) );
  CMXI2X1 U23557 ( .A0(n12986), .A1(n12980), .S(n4193), .Z(n12993) );
  CMX2X1 U23558 ( .A0(n12981), .A1(n12993), .S(n3810), .Z(n13010) );
  CMXI2X1 U23559 ( .A0(n12982), .A1(n13010), .S(n3469), .Z(N8455) );
  CMX2X1 U23560 ( .A0(N8089), .A1(N8088), .S(n3873), .Z(n12989) );
  CMXI2X1 U23561 ( .A0(n12989), .A1(n12983), .S(n4193), .Z(n13000) );
  CMX2X1 U23562 ( .A0(n12984), .A1(n13000), .S(n3811), .Z(n13013) );
  CMXI2X1 U23563 ( .A0(n12985), .A1(n13013), .S(n3468), .Z(N8456) );
  CMX2X1 U23564 ( .A0(N8088), .A1(N8087), .S(n3874), .Z(n12992) );
  CMX2X1 U23565 ( .A0(n12987), .A1(n13003), .S(n3812), .Z(n13016) );
  CMXI2X1 U23566 ( .A0(n12988), .A1(n13016), .S(n3467), .Z(N8457) );
  CMX2X1 U23567 ( .A0(N8087), .A1(N8086), .S(n3866), .Z(n12999) );
  CMXI2X1 U23568 ( .A0(n12999), .A1(n12989), .S(n4193), .Z(n13006) );
  CMX2X1 U23569 ( .A0(n12990), .A1(n13006), .S(n4369), .Z(n13019) );
  CMXI2X1 U23570 ( .A0(n12991), .A1(n13019), .S(n3466), .Z(N8458) );
  CMX2X1 U23571 ( .A0(N8086), .A1(N8085), .S(n3877), .Z(n13002) );
  CMXI2X1 U23572 ( .A0(n13002), .A1(n12992), .S(n4193), .Z(n13009) );
  CMX2X1 U23573 ( .A0(n12993), .A1(n13009), .S(n3771), .Z(n13022) );
  CMXI2X1 U23574 ( .A0(n12994), .A1(n13022), .S(n3465), .Z(N8459) );
  CMX2X1 U23575 ( .A0(n12996), .A1(n12995), .S(n3772), .Z(n15729) );
  CMX2X1 U23576 ( .A0(N8248), .A1(N8247), .S(n3869), .Z(n13062) );
  CMXI2X1 U23577 ( .A0(n13062), .A1(n12997), .S(n4193), .Z(n13134) );
  CMX2X1 U23578 ( .A0(n12998), .A1(n13134), .S(n3773), .Z(n13267) );
  CMXI2X1 U23579 ( .A0(n15729), .A1(n13267), .S(n3464), .Z(N8297) );
  CMX2X1 U23580 ( .A0(N8085), .A1(N8084), .S(n3870), .Z(n13005) );
  CMXI2X1 U23581 ( .A0(n13005), .A1(n12999), .S(n4193), .Z(n13012) );
  CMX2X1 U23582 ( .A0(n13000), .A1(n13012), .S(n3774), .Z(n13025) );
  CMXI2X1 U23583 ( .A0(n13001), .A1(n13025), .S(n3463), .Z(N8460) );
  CMX2X1 U23584 ( .A0(N8084), .A1(N8083), .S(n3871), .Z(n13008) );
  CMXI2X1 U23585 ( .A0(n13008), .A1(n13002), .S(n4193), .Z(n13015) );
  CMX2X1 U23586 ( .A0(n13003), .A1(n13015), .S(n3775), .Z(n13028) );
  CMXI2X1 U23587 ( .A0(n13004), .A1(n13028), .S(n3507), .Z(N8461) );
  CMX2X1 U23588 ( .A0(N8083), .A1(N8082), .S(n3872), .Z(n13011) );
  CMXI2X1 U23589 ( .A0(n13011), .A1(n13005), .S(n4193), .Z(n13018) );
  CMX2X1 U23590 ( .A0(n13006), .A1(n13018), .S(n3776), .Z(n13034) );
  CMXI2X1 U23591 ( .A0(n13007), .A1(n13034), .S(n3499), .Z(N8462) );
  CMX2X1 U23592 ( .A0(N8082), .A1(N8081), .S(n3873), .Z(n13014) );
  CMXI2X1 U23593 ( .A0(n13014), .A1(n13008), .S(n4193), .Z(n13021) );
  CMX2X1 U23594 ( .A0(n13009), .A1(n13021), .S(n3777), .Z(n13037) );
  CMXI2X1 U23595 ( .A0(n13010), .A1(n13037), .S(n3290), .Z(N8463) );
  CMX2X1 U23596 ( .A0(N8081), .A1(N8080), .S(n3874), .Z(n13017) );
  CMXI2X1 U23597 ( .A0(n13017), .A1(n13011), .S(n4193), .Z(n13024) );
  CMX2X1 U23598 ( .A0(n13012), .A1(n13024), .S(n3790), .Z(n13040) );
  CMXI2X1 U23599 ( .A0(n13013), .A1(n13040), .S(n3290), .Z(N8464) );
  CMX2X1 U23600 ( .A0(N8080), .A1(N8079), .S(n3875), .Z(n13020) );
  CMXI2X1 U23601 ( .A0(n13020), .A1(n13014), .S(n4193), .Z(n13027) );
  CMX2X1 U23602 ( .A0(n13015), .A1(n13027), .S(n3791), .Z(n13043) );
  CMXI2X1 U23603 ( .A0(n13016), .A1(n13043), .S(n3290), .Z(N8465) );
  CMX2X1 U23604 ( .A0(N8079), .A1(N8078), .S(n3862), .Z(n13023) );
  CMXI2X1 U23605 ( .A0(n13023), .A1(n13017), .S(n4193), .Z(n13033) );
  CMX2X1 U23606 ( .A0(n13018), .A1(n13033), .S(n3797), .Z(n13046) );
  CMXI2X1 U23607 ( .A0(n13019), .A1(n13046), .S(n3290), .Z(N8466) );
  CMX2X1 U23608 ( .A0(N8078), .A1(N8077), .S(n3863), .Z(n13026) );
  CMXI2X1 U23609 ( .A0(n13026), .A1(n13020), .S(n4193), .Z(n13036) );
  CMX2X1 U23610 ( .A0(n13021), .A1(n13036), .S(n3777), .Z(n13049) );
  CMXI2X1 U23611 ( .A0(n13022), .A1(n13049), .S(n3290), .Z(N8467) );
  CMX2X1 U23612 ( .A0(N8077), .A1(N8076), .S(n3876), .Z(n13032) );
  CMXI2X1 U23613 ( .A0(n13032), .A1(n13023), .S(n4193), .Z(n13039) );
  CMX2X1 U23614 ( .A0(n13024), .A1(n13039), .S(n3805), .Z(n13052) );
  CMXI2X1 U23615 ( .A0(n13025), .A1(n13052), .S(n3290), .Z(N8468) );
  CMX2X1 U23616 ( .A0(N8076), .A1(N8075), .S(n3877), .Z(n13035) );
  CMXI2X1 U23617 ( .A0(n13035), .A1(n13026), .S(n4192), .Z(n13042) );
  CMX2X1 U23618 ( .A0(n13027), .A1(n13042), .S(n3806), .Z(n13055) );
  CMXI2X1 U23619 ( .A0(n13028), .A1(n13055), .S(n3290), .Z(N8469) );
  CMX2X1 U23620 ( .A0(N8247), .A1(N8246), .S(n3869), .Z(n13100) );
  CMXI2X1 U23621 ( .A0(n13100), .A1(n13029), .S(n4192), .Z(n13167) );
  CMX2X1 U23622 ( .A0(n13030), .A1(n13167), .S(n3807), .Z(n13300) );
  CMXI2X1 U23623 ( .A0(n13031), .A1(n13300), .S(n3290), .Z(N8298) );
  CMX2X1 U23624 ( .A0(N8075), .A1(N8074), .S(n3870), .Z(n13038) );
  CMXI2X1 U23625 ( .A0(n13038), .A1(n13032), .S(n4192), .Z(n13045) );
  CMX2X1 U23626 ( .A0(n13033), .A1(n13045), .S(n3808), .Z(n13058) );
  CMX2X1 U23627 ( .A0(N8074), .A1(N8073), .S(n3871), .Z(n13041) );
  CMXI2X1 U23628 ( .A0(n13041), .A1(n13035), .S(n4192), .Z(n13048) );
  CMX2X1 U23629 ( .A0(n13036), .A1(n13048), .S(n3809), .Z(n13061) );
  CMX2X1 U23630 ( .A0(N8073), .A1(N8072), .S(n3872), .Z(n13044) );
  CMXI2X1 U23631 ( .A0(n13044), .A1(n13038), .S(n4192), .Z(n13051) );
  CMX2X1 U23632 ( .A0(n13039), .A1(n13051), .S(n3811), .Z(n13072) );
  CMXI2X1 U23633 ( .A0(n13040), .A1(n13072), .S(n3292), .Z(N8472) );
  CMX2X1 U23634 ( .A0(N8072), .A1(N8071), .S(n3867), .Z(n13047) );
  CMXI2X1 U23635 ( .A0(n13047), .A1(n13041), .S(n4192), .Z(n13054) );
  CMX2X1 U23636 ( .A0(n13042), .A1(n13054), .S(n3792), .Z(n13075) );
  CMXI2X1 U23637 ( .A0(n13043), .A1(n13075), .S(n3292), .Z(N8473) );
  CMX2X1 U23638 ( .A0(N8071), .A1(N8070), .S(n3869), .Z(n13050) );
  CMXI2X1 U23639 ( .A0(n13050), .A1(n13044), .S(n4192), .Z(n13057) );
  CMX2X1 U23640 ( .A0(n13045), .A1(n13057), .S(n3793), .Z(n13078) );
  CMXI2X1 U23641 ( .A0(n13046), .A1(n13078), .S(n3292), .Z(N8474) );
  CMX2X1 U23642 ( .A0(N8070), .A1(N8069), .S(n3870), .Z(n13053) );
  CMXI2X1 U23643 ( .A0(n13053), .A1(n13047), .S(n4192), .Z(n13060) );
  CMX2X1 U23644 ( .A0(n13048), .A1(n13060), .S(n3794), .Z(n13081) );
  CMXI2X1 U23645 ( .A0(n13049), .A1(n13081), .S(n3292), .Z(N8475) );
  CMX2X1 U23646 ( .A0(N8069), .A1(N8068), .S(n3878), .Z(n13056) );
  CMXI2X1 U23647 ( .A0(n13056), .A1(n13050), .S(n4192), .Z(n13071) );
  CMX2X1 U23648 ( .A0(n13051), .A1(n13071), .S(n3795), .Z(n13084) );
  CMXI2X1 U23649 ( .A0(n13052), .A1(n13084), .S(n3292), .Z(N8476) );
  CMX2X1 U23650 ( .A0(N8068), .A1(N8067), .S(n3878), .Z(n13059) );
  CMXI2X1 U23651 ( .A0(n13059), .A1(n13053), .S(n4192), .Z(n13074) );
  CMX2X1 U23652 ( .A0(n13054), .A1(n13074), .S(n3796), .Z(n13087) );
  CMXI2X1 U23653 ( .A0(n13055), .A1(n13087), .S(n3291), .Z(N8477) );
  CMX2X1 U23654 ( .A0(N8067), .A1(N8066), .S(n3879), .Z(n13070) );
  CMXI2X1 U23655 ( .A0(n13070), .A1(n13056), .S(n4192), .Z(n13077) );
  CMX2X1 U23656 ( .A0(n13057), .A1(n13077), .S(n3797), .Z(n13090) );
  CMXI2X1 U23657 ( .A0(n13058), .A1(n13090), .S(n3291), .Z(N8478) );
  CMX2X1 U23658 ( .A0(N8066), .A1(N8065), .S(n3880), .Z(n13073) );
  CMXI2X1 U23659 ( .A0(n13073), .A1(n13059), .S(n4192), .Z(n13080) );
  CMX2X1 U23660 ( .A0(n13060), .A1(n13080), .S(n3805), .Z(n13093) );
  CMXI2X1 U23661 ( .A0(n13061), .A1(n13093), .S(n3291), .Z(N8479) );
  CMX2X1 U23662 ( .A0(N8246), .A1(N8245), .S(n3881), .Z(n13133) );
  CMXI2X1 U23663 ( .A0(n13133), .A1(n13062), .S(n4192), .Z(n13200) );
  CMX2X1 U23664 ( .A0(n13063), .A1(n13200), .S(n3806), .Z(n13333) );
  CMXI2X1 U23665 ( .A0(n13064), .A1(n13333), .S(n3291), .Z(N8299) );
  CMXI2X1 U23666 ( .A0(n13737), .A1(n13740), .S(n4192), .Z(n14408) );
  CMXI2X1 U23667 ( .A0(N8276), .A1(N8275), .S(n3878), .Z(n13739) );
  CMXI2X1 U23668 ( .A0(N8277), .A1(N8278), .S(n3889), .Z(n13065) );
  CMXI2X1 U23669 ( .A0(n13739), .A1(n13065), .S(n4192), .Z(n13066) );
  CMXI2X1 U23670 ( .A0(n14408), .A1(n13066), .S(n3781), .Z(n13069) );
  CMXI2X1 U23671 ( .A0(N8269), .A1(N8270), .S(n3882), .Z(n13738) );
  CMXI2X1 U23672 ( .A0(n13067), .A1(n4433), .S(n4192), .Z(n14407) );
  CMX2X1 U23673 ( .A0(n14407), .A1(n13068), .S(n3807), .Z(n15730) );
  CMXI2X1 U23674 ( .A0(n13069), .A1(n15730), .S(n3291), .Z(N8281) );
  CMX2X1 U23675 ( .A0(N8065), .A1(N8064), .S(n3862), .Z(n13076) );
  CMXI2X1 U23676 ( .A0(n13076), .A1(n13070), .S(n4191), .Z(n13083) );
  CMX2X1 U23677 ( .A0(n13071), .A1(n13083), .S(n3808), .Z(n13096) );
  CMXI2X1 U23678 ( .A0(n13072), .A1(n13096), .S(n3291), .Z(N8480) );
  CMX2X1 U23679 ( .A0(N8064), .A1(N8063), .S(n3863), .Z(n13079) );
  CMXI2X1 U23680 ( .A0(n13079), .A1(n13073), .S(n4191), .Z(n13086) );
  CMX2X1 U23681 ( .A0(n13074), .A1(n13086), .S(n3809), .Z(n13099) );
  CMXI2X1 U23682 ( .A0(n13075), .A1(n13099), .S(n3291), .Z(N8481) );
  CMX2X1 U23683 ( .A0(N8063), .A1(N8062), .S(n3864), .Z(n13082) );
  CMXI2X1 U23684 ( .A0(n13082), .A1(n13076), .S(n4191), .Z(n13089) );
  CMX2X1 U23685 ( .A0(n13077), .A1(n13089), .S(n3810), .Z(n13105) );
  CMXI2X1 U23686 ( .A0(n13078), .A1(n13105), .S(n3291), .Z(N8482) );
  CMX2X1 U23687 ( .A0(N8062), .A1(N8061), .S(n3864), .Z(n13085) );
  CMXI2X1 U23688 ( .A0(n13085), .A1(n13079), .S(n4191), .Z(n13092) );
  CMX2X1 U23689 ( .A0(n13080), .A1(n13092), .S(n3811), .Z(n13108) );
  CMXI2X1 U23690 ( .A0(n13081), .A1(n13108), .S(n3291), .Z(N8483) );
  CMX2X1 U23691 ( .A0(N8061), .A1(N8060), .S(n3865), .Z(n13088) );
  CMXI2X1 U23692 ( .A0(n13088), .A1(n13082), .S(n4191), .Z(n13095) );
  CMX2X1 U23693 ( .A0(n13083), .A1(n13095), .S(n3812), .Z(n13111) );
  CMXI2X1 U23694 ( .A0(n13084), .A1(n13111), .S(n3291), .Z(N8484) );
  CMX2X1 U23695 ( .A0(N8060), .A1(N8059), .S(n3865), .Z(n13091) );
  CMXI2X1 U23696 ( .A0(n13091), .A1(n13085), .S(n4191), .Z(n13098) );
  CMX2X1 U23697 ( .A0(n13086), .A1(n13098), .S(n4366), .Z(n13114) );
  CMXI2X1 U23698 ( .A0(n13087), .A1(n13114), .S(n3291), .Z(N8485) );
  CMX2X1 U23699 ( .A0(N8059), .A1(N8058), .S(n3866), .Z(n13094) );
  CMXI2X1 U23700 ( .A0(n13094), .A1(n13088), .S(n4191), .Z(n13104) );
  CMX2X1 U23701 ( .A0(n13089), .A1(n13104), .S(n3771), .Z(n13117) );
  CMXI2X1 U23702 ( .A0(n13090), .A1(n13117), .S(n3294), .Z(N8486) );
  CMX2X1 U23703 ( .A0(N8058), .A1(N8057), .S(n3873), .Z(n13097) );
  CMXI2X1 U23704 ( .A0(n13097), .A1(n13091), .S(n4191), .Z(n13107) );
  CMX2X1 U23705 ( .A0(n13092), .A1(n13107), .S(n3805), .Z(n13120) );
  CMXI2X1 U23706 ( .A0(n13093), .A1(n13120), .S(n3293), .Z(N8487) );
  CMX2X1 U23707 ( .A0(N8057), .A1(N8056), .S(n3874), .Z(n13103) );
  CMXI2X1 U23708 ( .A0(n13103), .A1(n13094), .S(n4191), .Z(n13110) );
  CMX2X1 U23709 ( .A0(n13095), .A1(n13110), .S(n3792), .Z(n13123) );
  CMXI2X1 U23710 ( .A0(n13096), .A1(n13123), .S(n3293), .Z(N8488) );
  CMX2X1 U23711 ( .A0(N8056), .A1(N8055), .S(n3875), .Z(n13106) );
  CMXI2X1 U23712 ( .A0(n13106), .A1(n13097), .S(n4191), .Z(n13113) );
  CMX2X1 U23713 ( .A0(n13098), .A1(n13113), .S(n3772), .Z(n13126) );
  CMXI2X1 U23714 ( .A0(n13099), .A1(n13126), .S(n3293), .Z(N8489) );
  CMX2X1 U23715 ( .A0(N8245), .A1(N8244), .S(n3876), .Z(n13166) );
  CMXI2X1 U23716 ( .A0(n13166), .A1(n13100), .S(n4191), .Z(n13233) );
  CMX2X1 U23717 ( .A0(n13101), .A1(n13233), .S(n3773), .Z(n13366) );
  CMXI2X1 U23718 ( .A0(n13102), .A1(n13366), .S(n3293), .Z(N8300) );
  CMX2X1 U23719 ( .A0(N8055), .A1(N8054), .S(n3871), .Z(n13109) );
  CMXI2X1 U23720 ( .A0(n13109), .A1(n13103), .S(n4191), .Z(n13116) );
  CMX2X1 U23721 ( .A0(n13104), .A1(n13116), .S(n3774), .Z(n13129) );
  CMXI2X1 U23722 ( .A0(n13105), .A1(n13129), .S(n3293), .Z(N8490) );
  CMX2X1 U23723 ( .A0(N8054), .A1(N8053), .S(n3872), .Z(n13112) );
  CMXI2X1 U23724 ( .A0(n13112), .A1(n13106), .S(n4191), .Z(n13119) );
  CMX2X1 U23725 ( .A0(n13107), .A1(n13119), .S(n3775), .Z(n13132) );
  CMXI2X1 U23726 ( .A0(n13108), .A1(n13132), .S(n3293), .Z(N8491) );
  CMX2X1 U23727 ( .A0(N8053), .A1(N8052), .S(n3873), .Z(n13115) );
  CMXI2X1 U23728 ( .A0(n13115), .A1(n13109), .S(n4191), .Z(n13122) );
  CMX2X1 U23729 ( .A0(n13110), .A1(n13122), .S(n3776), .Z(n13138) );
  CMXI2X1 U23730 ( .A0(n13111), .A1(n13138), .S(n3293), .Z(N8492) );
  CMX2X1 U23731 ( .A0(N8052), .A1(N8051), .S(n3874), .Z(n13118) );
  CMXI2X1 U23732 ( .A0(n13118), .A1(n13112), .S(n4191), .Z(n13125) );
  CMX2X1 U23733 ( .A0(n13113), .A1(n13125), .S(n3777), .Z(n13141) );
  CMXI2X1 U23734 ( .A0(n13114), .A1(n13141), .S(n3293), .Z(N8493) );
  CMX2X1 U23735 ( .A0(N8051), .A1(N8050), .S(n3879), .Z(n13121) );
  CMXI2X1 U23736 ( .A0(n13121), .A1(n13115), .S(n4191), .Z(n13128) );
  CMX2X1 U23737 ( .A0(n13116), .A1(n13128), .S(n3790), .Z(n13144) );
  CMXI2X1 U23738 ( .A0(n13117), .A1(n13144), .S(n3293), .Z(N8494) );
  CMX2X1 U23739 ( .A0(N8050), .A1(N8049), .S(n3867), .Z(n13124) );
  CMXI2X1 U23740 ( .A0(n13124), .A1(n13118), .S(n4190), .Z(n13131) );
  CMX2X1 U23741 ( .A0(n13119), .A1(n13131), .S(n3791), .Z(n13147) );
  CMXI2X1 U23742 ( .A0(n13120), .A1(n13147), .S(n3293), .Z(N8495) );
  CMX2X1 U23743 ( .A0(N8049), .A1(N8048), .S(n3868), .Z(n13127) );
  CMXI2X1 U23744 ( .A0(n13127), .A1(n13121), .S(n4190), .Z(n13137) );
  CMX2X1 U23745 ( .A0(n13122), .A1(n13137), .S(n3792), .Z(n13150) );
  CMXI2X1 U23746 ( .A0(n13123), .A1(n13150), .S(n3293), .Z(N8496) );
  CMX2X1 U23747 ( .A0(N8048), .A1(N8047), .S(n3869), .Z(n13130) );
  CMXI2X1 U23748 ( .A0(n13130), .A1(n13124), .S(n4190), .Z(n13140) );
  CMX2X1 U23749 ( .A0(n13125), .A1(n13140), .S(n3793), .Z(n13153) );
  CMXI2X1 U23750 ( .A0(n13126), .A1(n13153), .S(n3292), .Z(N8497) );
  CMX2X1 U23751 ( .A0(N8047), .A1(N8046), .S(n3870), .Z(n13136) );
  CMXI2X1 U23752 ( .A0(n13136), .A1(n13127), .S(n4190), .Z(n13143) );
  CMX2X1 U23753 ( .A0(n13128), .A1(n13143), .S(n3794), .Z(n13156) );
  CMXI2X1 U23754 ( .A0(n13129), .A1(n13156), .S(n3292), .Z(N8498) );
  CMX2X1 U23755 ( .A0(N8046), .A1(N8045), .S(n3871), .Z(n13139) );
  CMXI2X1 U23756 ( .A0(n13139), .A1(n13130), .S(n4190), .Z(n13146) );
  CMX2X1 U23757 ( .A0(n13131), .A1(n13146), .S(n3795), .Z(n13159) );
  CMXI2X1 U23758 ( .A0(n13132), .A1(n13159), .S(n3292), .Z(N8499) );
  CMX2X1 U23759 ( .A0(N8244), .A1(N8243), .S(n3872), .Z(n13199) );
  CMXI2X1 U23760 ( .A0(n13199), .A1(n13133), .S(n4190), .Z(n13266) );
  CMX2X1 U23761 ( .A0(n13134), .A1(n13266), .S(n3796), .Z(n13399) );
  CMXI2X1 U23762 ( .A0(n13135), .A1(n13399), .S(n3292), .Z(N8301) );
  CMX2X1 U23763 ( .A0(N8045), .A1(N8044), .S(n3873), .Z(n13142) );
  CMXI2X1 U23764 ( .A0(n13142), .A1(n13136), .S(n4190), .Z(n13149) );
  CMX2X1 U23765 ( .A0(n13137), .A1(n13149), .S(n3797), .Z(n13162) );
  CMXI2X1 U23766 ( .A0(n13138), .A1(n13162), .S(n3292), .Z(N8500) );
  CMX2X1 U23767 ( .A0(N8044), .A1(N8043), .S(n3866), .Z(n13145) );
  CMXI2X1 U23768 ( .A0(n13145), .A1(n13139), .S(n4190), .Z(n13152) );
  CMX2X1 U23769 ( .A0(n13140), .A1(n13152), .S(n3805), .Z(n13165) );
  CMXI2X1 U23770 ( .A0(n13141), .A1(n13165), .S(n3295), .Z(N8501) );
  CMX2X1 U23771 ( .A0(N8043), .A1(N8042), .S(n3867), .Z(n13148) );
  CMXI2X1 U23772 ( .A0(n13148), .A1(n13142), .S(n4190), .Z(n13155) );
  CMX2X1 U23773 ( .A0(n13143), .A1(n13155), .S(n3806), .Z(n13171) );
  CMXI2X1 U23774 ( .A0(n13144), .A1(n13171), .S(n3295), .Z(N8502) );
  CMX2X1 U23775 ( .A0(N8042), .A1(N8041), .S(n3874), .Z(n13151) );
  CMXI2X1 U23776 ( .A0(n13151), .A1(n13145), .S(n4190), .Z(n13158) );
  CMX2X1 U23777 ( .A0(n13146), .A1(n13158), .S(n3796), .Z(n13174) );
  CMXI2X1 U23778 ( .A0(n13147), .A1(n13174), .S(n3295), .Z(N8503) );
  CMX2X1 U23779 ( .A0(N8041), .A1(N8040), .S(n3875), .Z(n13154) );
  CMXI2X1 U23780 ( .A0(n13154), .A1(n13148), .S(n4190), .Z(n13161) );
  CMX2X1 U23781 ( .A0(n13149), .A1(n13161), .S(n3773), .Z(n13177) );
  CMXI2X1 U23782 ( .A0(n13150), .A1(n13177), .S(n3295), .Z(N8504) );
  CMX2X1 U23783 ( .A0(N8040), .A1(N8039), .S(n3877), .Z(n13157) );
  CMXI2X1 U23784 ( .A0(n13157), .A1(n13151), .S(n4190), .Z(n13164) );
  CMX2X1 U23785 ( .A0(n13152), .A1(n13164), .S(n3811), .Z(n13180) );
  CMXI2X1 U23786 ( .A0(n13153), .A1(n13180), .S(n3295), .Z(N8505) );
  CMX2X1 U23787 ( .A0(N8039), .A1(N8038), .S(n3878), .Z(n13160) );
  CMXI2X1 U23788 ( .A0(n13160), .A1(n13154), .S(n4190), .Z(n13170) );
  CMX2X1 U23789 ( .A0(n13155), .A1(n13170), .S(n3812), .Z(n13183) );
  CMXI2X1 U23790 ( .A0(n13156), .A1(n13183), .S(n3295), .Z(N8506) );
  CMX2X1 U23791 ( .A0(N8038), .A1(N8037), .S(n3879), .Z(n13163) );
  CMXI2X1 U23792 ( .A0(n13163), .A1(n13157), .S(n4190), .Z(n13173) );
  CMX2X1 U23793 ( .A0(n13158), .A1(n13173), .S(n3771), .Z(n13186) );
  CMXI2X1 U23794 ( .A0(n13159), .A1(n13186), .S(n3295), .Z(N8507) );
  CMX2X1 U23795 ( .A0(N8037), .A1(N8036), .S(n3880), .Z(n13169) );
  CMXI2X1 U23796 ( .A0(n13169), .A1(n13160), .S(n4190), .Z(n13176) );
  CMX2X1 U23797 ( .A0(n13161), .A1(n13176), .S(n3792), .Z(n13189) );
  CMXI2X1 U23798 ( .A0(n13162), .A1(n13189), .S(n3295), .Z(N8508) );
  CMXI2X1 U23799 ( .A0(n13172), .A1(n13163), .S(n4190), .Z(n13179) );
  CMX2X1 U23800 ( .A0(n13164), .A1(n13179), .S(n3793), .Z(n13192) );
  CMXI2X1 U23801 ( .A0(n13165), .A1(n13192), .S(n3294), .Z(N8509) );
  CMX2X1 U23802 ( .A0(N8243), .A1(N8242), .S(n3876), .Z(n13232) );
  CMXI2X1 U23803 ( .A0(n13232), .A1(n13166), .S(n4189), .Z(n13299) );
  CMX2X1 U23804 ( .A0(n13167), .A1(n13299), .S(n3794), .Z(n13439) );
  CMXI2X1 U23805 ( .A0(n13168), .A1(n13439), .S(n3294), .Z(N8302) );
  CMX2X1 U23806 ( .A0(N8035), .A1(N8034), .S(n3877), .Z(n13175) );
  CMX2X1 U23807 ( .A0(n13170), .A1(n13182), .S(n3795), .Z(n13195) );
  CMXI2X1 U23808 ( .A0(n13171), .A1(n13195), .S(n3294), .Z(N8510) );
  CMX2X1 U23809 ( .A0(N8034), .A1(N8033), .S(n3878), .Z(n13178) );
  CMX2X1 U23810 ( .A0(n13173), .A1(n13185), .S(n3796), .Z(n13198) );
  CMXI2X1 U23811 ( .A0(n13174), .A1(n13198), .S(n3294), .Z(N8511) );
  CMX2X1 U23812 ( .A0(N8033), .A1(N8032), .S(n3880), .Z(n13181) );
  CMXI2X1 U23813 ( .A0(n13181), .A1(n13175), .S(n4189), .Z(n13188) );
  CMX2X1 U23814 ( .A0(n13176), .A1(n13188), .S(n3805), .Z(n13204) );
  CMXI2X1 U23815 ( .A0(n13177), .A1(n13204), .S(n3294), .Z(N8512) );
  CMX2X1 U23816 ( .A0(N8032), .A1(N8031), .S(n3876), .Z(n13184) );
  CMXI2X1 U23817 ( .A0(n13184), .A1(n13178), .S(n4189), .Z(n13191) );
  CMX2X1 U23818 ( .A0(n13179), .A1(n13191), .S(n3792), .Z(n13207) );
  CMXI2X1 U23819 ( .A0(n13180), .A1(n13207), .S(n3294), .Z(N8513) );
  CMX2X1 U23820 ( .A0(N8031), .A1(N8030), .S(n3877), .Z(n13187) );
  CMX2X1 U23821 ( .A0(n13182), .A1(n13194), .S(n3793), .Z(n13210) );
  CMXI2X1 U23822 ( .A0(n13183), .A1(n13210), .S(n3294), .Z(N8514) );
  CMX2X1 U23823 ( .A0(N8030), .A1(N8029), .S(n3878), .Z(n13190) );
  CMXI2X1 U23824 ( .A0(n13190), .A1(n13184), .S(n4189), .Z(n13197) );
  CMX2X1 U23825 ( .A0(n13185), .A1(n13197), .S(n3794), .Z(n13213) );
  CMXI2X1 U23826 ( .A0(n13186), .A1(n13213), .S(n3294), .Z(N8515) );
  CMX2X1 U23827 ( .A0(N8029), .A1(N8028), .S(n3879), .Z(n13193) );
  CMXI2X1 U23828 ( .A0(n13193), .A1(n13187), .S(n4189), .Z(n13203) );
  CMX2X1 U23829 ( .A0(n13188), .A1(n13203), .S(n3795), .Z(n13216) );
  CMXI2X1 U23830 ( .A0(n13189), .A1(n13216), .S(n3294), .Z(N8516) );
  CMX2X1 U23831 ( .A0(N8028), .A1(N8027), .S(n3880), .Z(n13196) );
  CMXI2X1 U23832 ( .A0(n13196), .A1(n13190), .S(n4189), .Z(n13206) );
  CMX2X1 U23833 ( .A0(n13191), .A1(n13206), .S(n3796), .Z(n13219) );
  CMXI2X1 U23834 ( .A0(n13192), .A1(n13219), .S(n3294), .Z(N8517) );
  CMX2X1 U23835 ( .A0(N8027), .A1(N8026), .S(n3881), .Z(n13202) );
  CMXI2X1 U23836 ( .A0(n13202), .A1(n13193), .S(n4189), .Z(n13209) );
  CMX2X1 U23837 ( .A0(n13194), .A1(n13209), .S(n3797), .Z(n13222) );
  CMXI2X1 U23838 ( .A0(n13195), .A1(n13222), .S(n3297), .Z(N8518) );
  CMX2X1 U23839 ( .A0(N8026), .A1(N8025), .S(n3862), .Z(n13205) );
  CMXI2X1 U23840 ( .A0(n13205), .A1(n13196), .S(n4189), .Z(n13212) );
  CMX2X1 U23841 ( .A0(n13197), .A1(n13212), .S(n3805), .Z(n13225) );
  CMXI2X1 U23842 ( .A0(n13198), .A1(n13225), .S(n3297), .Z(N8519) );
  CMX2X1 U23843 ( .A0(N8242), .A1(N8241), .S(n3868), .Z(n13265) );
  CMXI2X1 U23844 ( .A0(n13265), .A1(n13199), .S(n4189), .Z(n13332) );
  CMX2X1 U23845 ( .A0(n13200), .A1(n13332), .S(n3806), .Z(n13472) );
  CMXI2X1 U23846 ( .A0(n13201), .A1(n13472), .S(n3297), .Z(N8303) );
  CMX2X1 U23847 ( .A0(N8025), .A1(N8024), .S(n3869), .Z(n13208) );
  CMXI2X1 U23848 ( .A0(n13208), .A1(n13202), .S(n4189), .Z(n13215) );
  CMX2X1 U23849 ( .A0(n13203), .A1(n13215), .S(n3807), .Z(n13228) );
  CMXI2X1 U23850 ( .A0(n13204), .A1(n13228), .S(n3296), .Z(N8520) );
  CMX2X1 U23851 ( .A0(N8024), .A1(N8023), .S(n3863), .Z(n13211) );
  CMXI2X1 U23852 ( .A0(n13211), .A1(n13205), .S(n4189), .Z(n13218) );
  CMX2X1 U23853 ( .A0(n13206), .A1(n13218), .S(n3808), .Z(n13231) );
  CMXI2X1 U23854 ( .A0(n13207), .A1(n13231), .S(n3296), .Z(N8521) );
  CMX2X1 U23855 ( .A0(N8023), .A1(N8022), .S(n3864), .Z(n13214) );
  CMXI2X1 U23856 ( .A0(n13214), .A1(n13208), .S(n4189), .Z(n13221) );
  CMX2X1 U23857 ( .A0(n13209), .A1(n13221), .S(n3809), .Z(n13237) );
  CMXI2X1 U23858 ( .A0(n13210), .A1(n13237), .S(n3296), .Z(N8522) );
  CMX2X1 U23859 ( .A0(N8022), .A1(N8021), .S(n3881), .Z(n13217) );
  CMXI2X1 U23860 ( .A0(n13217), .A1(n13211), .S(n4189), .Z(n13224) );
  CMX2X1 U23861 ( .A0(n13212), .A1(n13224), .S(n3810), .Z(n13240) );
  CMXI2X1 U23862 ( .A0(n13213), .A1(n13240), .S(n3296), .Z(N8523) );
  CMX2X1 U23863 ( .A0(N8021), .A1(N8020), .S(n3862), .Z(n13220) );
  CMXI2X1 U23864 ( .A0(n13220), .A1(n13214), .S(n4188), .Z(n13227) );
  CMX2X1 U23865 ( .A0(n13215), .A1(n13227), .S(n3811), .Z(n13243) );
  CMXI2X1 U23866 ( .A0(n13216), .A1(n13243), .S(n3296), .Z(N8524) );
  CMX2X1 U23867 ( .A0(N8020), .A1(N8019), .S(n3863), .Z(n13223) );
  CMXI2X1 U23868 ( .A0(n13223), .A1(n13217), .S(n4188), .Z(n13230) );
  CMX2X1 U23869 ( .A0(n13218), .A1(n13230), .S(n3812), .Z(n13246) );
  CMX2X1 U23870 ( .A0(N8019), .A1(N8018), .S(n3864), .Z(n13226) );
  CMXI2X1 U23871 ( .A0(n13226), .A1(n13220), .S(n4188), .Z(n13236) );
  CMX2X1 U23872 ( .A0(n13221), .A1(n13236), .S(n4373), .Z(n13249) );
  CMXI2X1 U23873 ( .A0(n13222), .A1(n13249), .S(n3296), .Z(N8526) );
  CMX2X1 U23874 ( .A0(N8018), .A1(N8017), .S(n3879), .Z(n13229) );
  CMXI2X1 U23875 ( .A0(n13229), .A1(n13223), .S(n4188), .Z(n13239) );
  CMX2X1 U23876 ( .A0(n13224), .A1(n13239), .S(n3771), .Z(n13252) );
  CMXI2X1 U23877 ( .A0(n13225), .A1(n13252), .S(n3296), .Z(N8527) );
  CMX2X1 U23878 ( .A0(N8017), .A1(N8016), .S(n3880), .Z(n13235) );
  CMX2X1 U23879 ( .A0(n13227), .A1(n13242), .S(n3792), .Z(n13255) );
  CMXI2X1 U23880 ( .A0(n13228), .A1(n13255), .S(n3296), .Z(N8528) );
  CMX2X1 U23881 ( .A0(N8016), .A1(N8015), .S(n3881), .Z(n13238) );
  CMXI2X1 U23882 ( .A0(n13238), .A1(n13229), .S(n4188), .Z(n13245) );
  CMX2X1 U23883 ( .A0(n13230), .A1(n13245), .S(n3772), .Z(n13258) );
  CMXI2X1 U23884 ( .A0(n13231), .A1(n13258), .S(n3296), .Z(N8529) );
  CMX2X1 U23885 ( .A0(N8241), .A1(N8240), .S(n3862), .Z(n13298) );
  CMXI2X1 U23886 ( .A0(n13298), .A1(n13232), .S(n4188), .Z(n13365) );
  CMX2X1 U23887 ( .A0(n13233), .A1(n13365), .S(n3797), .Z(n13505) );
  CMXI2X1 U23888 ( .A0(n13234), .A1(n13505), .S(n3296), .Z(N8304) );
  CMX2X1 U23889 ( .A0(N8015), .A1(N8014), .S(n3881), .Z(n13241) );
  CMXI2X1 U23890 ( .A0(n13241), .A1(n13235), .S(n4188), .Z(n13248) );
  CMX2X1 U23891 ( .A0(n13236), .A1(n13248), .S(n3805), .Z(n13261) );
  CMXI2X1 U23892 ( .A0(n13237), .A1(n13261), .S(n3296), .Z(N8530) );
  CMX2X1 U23893 ( .A0(N8014), .A1(N8013), .S(n3865), .Z(n13244) );
  CMXI2X1 U23894 ( .A0(n13244), .A1(n13238), .S(n4188), .Z(n13251) );
  CMX2X1 U23895 ( .A0(n13239), .A1(n13251), .S(n3806), .Z(n13264) );
  CMXI2X1 U23896 ( .A0(n13240), .A1(n13264), .S(n3295), .Z(N8531) );
  CMX2X1 U23897 ( .A0(N8013), .A1(N8012), .S(n3866), .Z(n13247) );
  CMXI2X1 U23898 ( .A0(n13247), .A1(n13241), .S(n4188), .Z(n13254) );
  CMX2X1 U23899 ( .A0(n13242), .A1(n13254), .S(n3807), .Z(n13270) );
  CMXI2X1 U23900 ( .A0(n13243), .A1(n13270), .S(n3295), .Z(N8532) );
  CMX2X1 U23901 ( .A0(N8012), .A1(N8011), .S(n3867), .Z(n13250) );
  CMXI2X1 U23902 ( .A0(n13250), .A1(n13244), .S(n4188), .Z(n13257) );
  CMX2X1 U23903 ( .A0(n13245), .A1(n13257), .S(n3808), .Z(n13273) );
  CMXI2X1 U23904 ( .A0(n13246), .A1(n13273), .S(n3295), .Z(N8533) );
  CMX2X1 U23905 ( .A0(N8011), .A1(N8010), .S(n3868), .Z(n13253) );
  CMXI2X1 U23906 ( .A0(n13253), .A1(n13247), .S(n4188), .Z(n13260) );
  CMX2X1 U23907 ( .A0(n13248), .A1(n13260), .S(n3806), .Z(n13276) );
  CMXI2X1 U23908 ( .A0(n13249), .A1(n13276), .S(n3298), .Z(N8534) );
  CMX2X1 U23909 ( .A0(N8010), .A1(N8009), .S(n3869), .Z(n13256) );
  CMXI2X1 U23910 ( .A0(n13256), .A1(n13250), .S(n4188), .Z(n13263) );
  CMX2X1 U23911 ( .A0(n13251), .A1(n13263), .S(n3772), .Z(n13279) );
  CMXI2X1 U23912 ( .A0(n13252), .A1(n13279), .S(n3298), .Z(N8535) );
  CMX2X1 U23913 ( .A0(N8009), .A1(N8008), .S(n3870), .Z(n13259) );
  CMXI2X1 U23914 ( .A0(n13259), .A1(n13253), .S(n4188), .Z(n13269) );
  CMX2X1 U23915 ( .A0(n13254), .A1(n13269), .S(n3773), .Z(n13282) );
  CMXI2X1 U23916 ( .A0(n13255), .A1(n13282), .S(n3298), .Z(N8536) );
  CMX2X1 U23917 ( .A0(N8008), .A1(N8007), .S(n3871), .Z(n13262) );
  CMXI2X1 U23918 ( .A0(n13262), .A1(n13256), .S(n4188), .Z(n13272) );
  CMX2X1 U23919 ( .A0(n13257), .A1(n13272), .S(n3774), .Z(n13285) );
  CMXI2X1 U23920 ( .A0(n13258), .A1(n13285), .S(n3298), .Z(N8537) );
  CMX2X1 U23921 ( .A0(N8007), .A1(N8006), .S(n3870), .Z(n13268) );
  CMXI2X1 U23922 ( .A0(n13268), .A1(n13259), .S(n4188), .Z(n13275) );
  CMX2X1 U23923 ( .A0(n13260), .A1(n13275), .S(n3775), .Z(n13288) );
  CMXI2X1 U23924 ( .A0(n13261), .A1(n13288), .S(n3298), .Z(N8538) );
  CMX2X1 U23925 ( .A0(N8006), .A1(N8005), .S(n3871), .Z(n13271) );
  CMX2X1 U23926 ( .A0(n13263), .A1(n13278), .S(n3776), .Z(n13291) );
  CMXI2X1 U23927 ( .A0(n13264), .A1(n13291), .S(n3298), .Z(N8539) );
  CMX2X1 U23928 ( .A0(N8240), .A1(N8239), .S(n3872), .Z(n13331) );
  CMXI2X1 U23929 ( .A0(n13331), .A1(n13265), .S(n4187), .Z(n13398) );
  CMX2X1 U23930 ( .A0(n13266), .A1(n13398), .S(n3777), .Z(n13538) );
  CMXI2X1 U23931 ( .A0(n13267), .A1(n13538), .S(n3298), .Z(N8305) );
  CMX2X1 U23932 ( .A0(N8005), .A1(N8004), .S(n3873), .Z(n13274) );
  CMXI2X1 U23933 ( .A0(n13274), .A1(n13268), .S(n4187), .Z(n13281) );
  CMX2X1 U23934 ( .A0(n13269), .A1(n13281), .S(n3790), .Z(n13294) );
  CMXI2X1 U23935 ( .A0(n13270), .A1(n13294), .S(n3298), .Z(N8540) );
  CMX2X1 U23936 ( .A0(N8004), .A1(N8003), .S(n3865), .Z(n13277) );
  CMXI2X1 U23937 ( .A0(n13277), .A1(n13271), .S(n4187), .Z(n13284) );
  CMX2X1 U23938 ( .A0(n13272), .A1(n13284), .S(n3791), .Z(n13297) );
  CMXI2X1 U23939 ( .A0(n13273), .A1(n13297), .S(n3298), .Z(N8541) );
  CMX2X1 U23940 ( .A0(N8003), .A1(N8002), .S(n3866), .Z(n13280) );
  CMXI2X1 U23941 ( .A0(n13280), .A1(n13274), .S(n4187), .Z(n13287) );
  CMX2X1 U23942 ( .A0(n13275), .A1(n13287), .S(n3792), .Z(n13303) );
  CMXI2X1 U23943 ( .A0(n13276), .A1(n13303), .S(n3297), .Z(N8542) );
  CMX2X1 U23944 ( .A0(N8002), .A1(N8001), .S(n3867), .Z(n13283) );
  CMXI2X1 U23945 ( .A0(n13283), .A1(n13277), .S(n4187), .Z(n13290) );
  CMX2X1 U23946 ( .A0(n13278), .A1(n13290), .S(n3793), .Z(n13306) );
  CMXI2X1 U23947 ( .A0(n13279), .A1(n13306), .S(n3297), .Z(N8543) );
  CMX2X1 U23948 ( .A0(N8001), .A1(N8000), .S(n3868), .Z(n13286) );
  CMXI2X1 U23949 ( .A0(n13286), .A1(n13280), .S(n4187), .Z(n13293) );
  CMX2X1 U23950 ( .A0(n13281), .A1(n13293), .S(n3794), .Z(n13309) );
  CMXI2X1 U23951 ( .A0(n13282), .A1(n13309), .S(n3297), .Z(N8544) );
  CMX2X1 U23952 ( .A0(N8000), .A1(N7999), .S(n3863), .Z(n13289) );
  CMXI2X1 U23953 ( .A0(n13289), .A1(n13283), .S(n4187), .Z(n13296) );
  CMX2X1 U23954 ( .A0(n13284), .A1(n13296), .S(n3795), .Z(n13312) );
  CMXI2X1 U23955 ( .A0(n13285), .A1(n13312), .S(n3297), .Z(N8545) );
  CMX2X1 U23956 ( .A0(N7999), .A1(N7998), .S(n3864), .Z(n13292) );
  CMXI2X1 U23957 ( .A0(n13292), .A1(n13286), .S(n4187), .Z(n13302) );
  CMX2X1 U23958 ( .A0(n13287), .A1(n13302), .S(n3796), .Z(n13315) );
  CMXI2X1 U23959 ( .A0(n13288), .A1(n13315), .S(n3297), .Z(N8546) );
  CMX2X1 U23960 ( .A0(N7998), .A1(N7997), .S(n3865), .Z(n13295) );
  CMXI2X1 U23961 ( .A0(n13295), .A1(n13289), .S(n4187), .Z(n13305) );
  CMX2X1 U23962 ( .A0(n13290), .A1(n13305), .S(n3797), .Z(n13318) );
  CMXI2X1 U23963 ( .A0(n13291), .A1(n13318), .S(n3297), .Z(N8547) );
  CMX2X1 U23964 ( .A0(N7997), .A1(N7996), .S(n3866), .Z(n13301) );
  CMXI2X1 U23965 ( .A0(n13301), .A1(n13292), .S(n4187), .Z(n13308) );
  CMX2X1 U23966 ( .A0(n13293), .A1(n13308), .S(n3805), .Z(n13321) );
  CMXI2X1 U23967 ( .A0(n13294), .A1(n13321), .S(n3297), .Z(N8548) );
  CMX2X1 U23968 ( .A0(N7996), .A1(N7995), .S(n3862), .Z(n13304) );
  CMXI2X1 U23969 ( .A0(n13304), .A1(n13295), .S(n4187), .Z(n13311) );
  CMX2X1 U23970 ( .A0(n13296), .A1(n13311), .S(n3806), .Z(n13324) );
  CMX2X1 U23971 ( .A0(N8239), .A1(N8238), .S(n3874), .Z(n13364) );
  CMXI2X1 U23972 ( .A0(n13364), .A1(n13298), .S(n4187), .Z(n13438) );
  CMX2X1 U23973 ( .A0(n13299), .A1(n13438), .S(n3793), .Z(n13571) );
  CMXI2X1 U23974 ( .A0(n13300), .A1(n13571), .S(n3297), .Z(N8306) );
  CMX2X1 U23975 ( .A0(N7995), .A1(N7994), .S(n3875), .Z(n13307) );
  CMXI2X1 U23976 ( .A0(n13307), .A1(n13301), .S(n4187), .Z(n13314) );
  CMX2X1 U23977 ( .A0(n13302), .A1(n13314), .S(n3773), .Z(n13327) );
  CMXI2X1 U23978 ( .A0(n13303), .A1(n13327), .S(n3276), .Z(N8550) );
  CMX2X1 U23979 ( .A0(N7994), .A1(N7993), .S(n3876), .Z(n13310) );
  CMXI2X1 U23980 ( .A0(n13310), .A1(n13304), .S(n4187), .Z(n13317) );
  CMX2X1 U23981 ( .A0(n13305), .A1(n13317), .S(n3809), .Z(n13330) );
  CMXI2X1 U23982 ( .A0(n13306), .A1(n13330), .S(n3276), .Z(N8551) );
  CMX2X1 U23983 ( .A0(N7993), .A1(N7992), .S(n3877), .Z(n13313) );
  CMXI2X1 U23984 ( .A0(n13313), .A1(n13307), .S(n4187), .Z(n13320) );
  CMX2X1 U23985 ( .A0(n13308), .A1(n13320), .S(n3810), .Z(n13336) );
  CMXI2X1 U23986 ( .A0(n13309), .A1(n13336), .S(n3276), .Z(N8552) );
  CMX2X1 U23987 ( .A0(N7992), .A1(N7991), .S(n3878), .Z(n13316) );
  CMXI2X1 U23988 ( .A0(n13316), .A1(n13310), .S(n4186), .Z(n13323) );
  CMX2X1 U23989 ( .A0(n13311), .A1(n13323), .S(n3811), .Z(n13339) );
  CMXI2X1 U23990 ( .A0(n13312), .A1(n13339), .S(n3276), .Z(N8553) );
  CMX2X1 U23991 ( .A0(N7991), .A1(N7990), .S(n3879), .Z(n13319) );
  CMXI2X1 U23992 ( .A0(n13319), .A1(n13313), .S(n4186), .Z(n13326) );
  CMX2X1 U23993 ( .A0(n13314), .A1(n13326), .S(n3812), .Z(n13342) );
  CMXI2X1 U23994 ( .A0(n13315), .A1(n13342), .S(n3277), .Z(N8554) );
  CMX2X1 U23995 ( .A0(N7990), .A1(N7989), .S(n3880), .Z(n13322) );
  CMX2X1 U23996 ( .A0(n13317), .A1(n13329), .S(n4305), .Z(n13345) );
  CMXI2X1 U23997 ( .A0(n13318), .A1(n13345), .S(n3277), .Z(N8555) );
  CMX2X1 U23998 ( .A0(N7989), .A1(N7988), .S(n3872), .Z(n13325) );
  CMXI2X1 U23999 ( .A0(n13325), .A1(n13319), .S(n4186), .Z(n13335) );
  CMX2X1 U24000 ( .A0(n13320), .A1(n13335), .S(n3807), .Z(n13348) );
  CMXI2X1 U24001 ( .A0(n13321), .A1(n13348), .S(n3277), .Z(N8556) );
  CMX2X1 U24002 ( .A0(N7988), .A1(N7987), .S(n3873), .Z(n13328) );
  CMXI2X1 U24003 ( .A0(n13328), .A1(n13322), .S(n4186), .Z(n13338) );
  CMX2X1 U24004 ( .A0(n13323), .A1(n13338), .S(n3807), .Z(n13351) );
  CMXI2X1 U24005 ( .A0(n13324), .A1(n13351), .S(n3277), .Z(N8557) );
  CMX2X1 U24006 ( .A0(N7987), .A1(N7986), .S(n3881), .Z(n13334) );
  CMXI2X1 U24007 ( .A0(n13334), .A1(n13325), .S(n4186), .Z(n13341) );
  CMX2X1 U24008 ( .A0(n13326), .A1(n13341), .S(n3808), .Z(n13354) );
  CMXI2X1 U24009 ( .A0(n13327), .A1(n13354), .S(n3277), .Z(N8558) );
  CMX2X1 U24010 ( .A0(N7986), .A1(N7985), .S(n3862), .Z(n13337) );
  CMX2X1 U24011 ( .A0(n13329), .A1(n13344), .S(n3809), .Z(n13357) );
  CMXI2X1 U24012 ( .A0(n13330), .A1(n13357), .S(n3277), .Z(N8559) );
  CMX2X1 U24013 ( .A0(N8238), .A1(N8237), .S(n3868), .Z(n13397) );
  CMXI2X1 U24014 ( .A0(n13397), .A1(n13331), .S(n4186), .Z(n13471) );
  CMX2X1 U24015 ( .A0(n13332), .A1(n13471), .S(n3810), .Z(n13604) );
  CMXI2X1 U24016 ( .A0(n13333), .A1(n13604), .S(n3277), .Z(N8307) );
  CMX2X1 U24017 ( .A0(N7985), .A1(N7984), .S(n3867), .Z(n13340) );
  CMX2X1 U24018 ( .A0(n13335), .A1(n13347), .S(n3811), .Z(n13360) );
  CMXI2X1 U24019 ( .A0(n13336), .A1(n13360), .S(n3277), .Z(N8560) );
  CMX2X1 U24020 ( .A0(N7984), .A1(N7983), .S(n3868), .Z(n13343) );
  CMX2X1 U24021 ( .A0(n13338), .A1(n13350), .S(n3812), .Z(n13363) );
  CMXI2X1 U24022 ( .A0(n13339), .A1(n13363), .S(n3277), .Z(N8561) );
  CMX2X1 U24023 ( .A0(N7983), .A1(N7982), .S(n3867), .Z(n13346) );
  CMXI2X1 U24024 ( .A0(n13346), .A1(n13340), .S(n4186), .Z(n13353) );
  CMX2X1 U24025 ( .A0(n13341), .A1(n13353), .S(n4371), .Z(n13369) );
  CMXI2X1 U24026 ( .A0(n13342), .A1(n13369), .S(n3480), .Z(N8562) );
  CMX2X1 U24027 ( .A0(N7982), .A1(N7981), .S(n3869), .Z(n13349) );
  CMXI2X1 U24028 ( .A0(n13349), .A1(n13343), .S(n4186), .Z(n13356) );
  CMX2X1 U24029 ( .A0(n13344), .A1(n13356), .S(n3771), .Z(n13372) );
  CMXI2X1 U24030 ( .A0(n13345), .A1(n13372), .S(n3481), .Z(N8563) );
  CMX2X1 U24031 ( .A0(N7981), .A1(N7980), .S(n3870), .Z(n13352) );
  CMXI2X1 U24032 ( .A0(n13352), .A1(n13346), .S(n4186), .Z(n13359) );
  CMX2X1 U24033 ( .A0(n13347), .A1(n3744), .S(n3772), .Z(n13375) );
  CMXI2X1 U24034 ( .A0(n13348), .A1(n13375), .S(n3478), .Z(N8564) );
  CMX2X1 U24035 ( .A0(N7980), .A1(N7979), .S(n3871), .Z(n13355) );
  CMXI2X1 U24036 ( .A0(n13355), .A1(n13349), .S(n4186), .Z(n13362) );
  CMX2X1 U24037 ( .A0(n13350), .A1(n13362), .S(n3773), .Z(n13378) );
  CMXI2X1 U24038 ( .A0(n13351), .A1(n13378), .S(n3298), .Z(N8565) );
  CMX2X1 U24039 ( .A0(N7979), .A1(N7978), .S(n3872), .Z(n13358) );
  CMXI2X1 U24040 ( .A0(n13358), .A1(n13352), .S(n4186), .Z(n13368) );
  CMX2X1 U24041 ( .A0(n13353), .A1(n13368), .S(n3774), .Z(n13381) );
  CMXI2X1 U24042 ( .A0(n13354), .A1(n13381), .S(n3298), .Z(N8566) );
  CMX2X1 U24043 ( .A0(N7978), .A1(N7977), .S(n3864), .Z(n13361) );
  CMXI2X1 U24044 ( .A0(n13361), .A1(n13355), .S(n4186), .Z(n13371) );
  CMX2X1 U24045 ( .A0(n13356), .A1(n13371), .S(n3775), .Z(n13384) );
  CMXI2X1 U24046 ( .A0(n13357), .A1(n13384), .S(n3275), .Z(N8567) );
  CMX2X1 U24047 ( .A0(N7977), .A1(N7976), .S(n3874), .Z(n13367) );
  CMX2X1 U24048 ( .A0(n13359), .A1(n13374), .S(n3776), .Z(n13387) );
  CMXI2X1 U24049 ( .A0(n13360), .A1(n13387), .S(n3275), .Z(N8568) );
  CMX2X1 U24050 ( .A0(N7976), .A1(N7975), .S(n3875), .Z(n13370) );
  CMX2X1 U24051 ( .A0(n13362), .A1(n13377), .S(n3777), .Z(n13390) );
  CMXI2X1 U24052 ( .A0(n13363), .A1(n13390), .S(n3275), .Z(N8569) );
  CMX2X1 U24053 ( .A0(N8237), .A1(N8236), .S(n3876), .Z(n13437) );
  CMXI2X1 U24054 ( .A0(n13437), .A1(n13364), .S(n4185), .Z(n13504) );
  CMX2X1 U24055 ( .A0(n13365), .A1(n13504), .S(n3790), .Z(n13637) );
  CMXI2X1 U24056 ( .A0(n13366), .A1(n13637), .S(n3275), .Z(N8308) );
  CMX2X1 U24057 ( .A0(N7975), .A1(N7974), .S(n3877), .Z(n13373) );
  CMXI2X1 U24058 ( .A0(n13373), .A1(n13367), .S(n4185), .Z(n13380) );
  CMX2X1 U24059 ( .A0(n13368), .A1(n13380), .S(n3791), .Z(n13393) );
  CMXI2X1 U24060 ( .A0(n13369), .A1(n13393), .S(n3275), .Z(N8570) );
  CMX2X1 U24061 ( .A0(N7974), .A1(N7973), .S(n3864), .Z(n13376) );
  CMX2X1 U24062 ( .A0(n13371), .A1(n13383), .S(n3794), .Z(n13396) );
  CMXI2X1 U24063 ( .A0(n13372), .A1(n13396), .S(n3275), .Z(N8571) );
  CMX2X1 U24064 ( .A0(N7973), .A1(N7972), .S(n3866), .Z(n13379) );
  CMXI2X1 U24065 ( .A0(n13379), .A1(n13373), .S(n4185), .Z(n13386) );
  CMX2X1 U24066 ( .A0(n13374), .A1(n13386), .S(n3774), .Z(n13409) );
  CMXI2X1 U24067 ( .A0(n13375), .A1(n13409), .S(n3275), .Z(N8572) );
  CMX2X1 U24068 ( .A0(N7972), .A1(N7971), .S(n3867), .Z(n13382) );
  CMXI2X1 U24069 ( .A0(n13382), .A1(n13376), .S(n4185), .Z(n13389) );
  CMX2X1 U24070 ( .A0(n13377), .A1(n13389), .S(n3810), .Z(n13412) );
  CMXI2X1 U24071 ( .A0(n13378), .A1(n13412), .S(n3275), .Z(N8573) );
  CMX2X1 U24072 ( .A0(N7971), .A1(N7970), .S(n3868), .Z(n13385) );
  CMXI2X1 U24073 ( .A0(n13385), .A1(n13379), .S(n4185), .Z(n13392) );
  CMX2X1 U24074 ( .A0(n13380), .A1(n13392), .S(n3771), .Z(n13415) );
  CMXI2X1 U24075 ( .A0(n13381), .A1(n13415), .S(n3275), .Z(N8574) );
  CMX2X1 U24076 ( .A0(N7970), .A1(N7969), .S(n3869), .Z(n13388) );
  CMXI2X1 U24077 ( .A0(n13388), .A1(n13382), .S(n4185), .Z(n13395) );
  CMX2X1 U24078 ( .A0(n13383), .A1(n13395), .S(n4307), .Z(n13418) );
  CMX2X1 U24079 ( .A0(N7969), .A1(N7968), .S(n3870), .Z(n13391) );
  CMXI2X1 U24080 ( .A0(n13391), .A1(n13385), .S(n4185), .Z(n13408) );
  CMX2X1 U24081 ( .A0(n13386), .A1(n13408), .S(n4307), .Z(n13421) );
  CMXI2X1 U24082 ( .A0(n13387), .A1(n13421), .S(n3275), .Z(N8576) );
  CMX2X1 U24083 ( .A0(N7968), .A1(N7967), .S(n3871), .Z(n13394) );
  CMXI2X1 U24084 ( .A0(n13394), .A1(n13388), .S(n4185), .Z(n13411) );
  CMX2X1 U24085 ( .A0(n13389), .A1(n13411), .S(n4322), .Z(n13424) );
  CMXI2X1 U24086 ( .A0(n13390), .A1(n13424), .S(n3276), .Z(N8577) );
  CMX2X1 U24087 ( .A0(N7967), .A1(N7966), .S(n3872), .Z(n13407) );
  CMXI2X1 U24088 ( .A0(n13407), .A1(n13391), .S(n4185), .Z(n13414) );
  CMX2X1 U24089 ( .A0(n13392), .A1(n13414), .S(n4307), .Z(n13427) );
  CMXI2X1 U24090 ( .A0(n13393), .A1(n13427), .S(n3276), .Z(N8578) );
  CMX2X1 U24091 ( .A0(N7966), .A1(N7965), .S(n3867), .Z(n13410) );
  CMX2X1 U24092 ( .A0(n13395), .A1(n13417), .S(n4307), .Z(n13430) );
  CMXI2X1 U24093 ( .A0(n13396), .A1(n13430), .S(n3276), .Z(N8579) );
  CMX2X1 U24094 ( .A0(N8236), .A1(N8235), .S(n3868), .Z(n13470) );
  CMXI2X1 U24095 ( .A0(n13470), .A1(n13397), .S(n4185), .Z(n13537) );
  CMX2X1 U24096 ( .A0(n13398), .A1(n13537), .S(n4307), .Z(n13670) );
  CMXI2X1 U24097 ( .A0(n13399), .A1(n13670), .S(n3276), .Z(N8309) );
  CMXI2X1 U24098 ( .A0(n13401), .A1(n13400), .S(n4185), .Z(n14742) );
  CMXI2X1 U24099 ( .A0(n13406), .A1(n13405), .S(n3276), .Z(N8282) );
  CMX2X1 U24100 ( .A0(N7965), .A1(N7964), .S(n3873), .Z(n13413) );
  CMX2X1 U24101 ( .A0(n13408), .A1(n13420), .S(n4307), .Z(n13433) );
  CMXI2X1 U24102 ( .A0(n13409), .A1(n13433), .S(n3276), .Z(N8580) );
  CMX2X1 U24103 ( .A0(N7964), .A1(N7963), .S(n3874), .Z(n13416) );
  CMXI2X1 U24104 ( .A0(n13416), .A1(n13410), .S(n4184), .Z(n13423) );
  CMX2X1 U24105 ( .A0(n13411), .A1(n13423), .S(n4307), .Z(n13436) );
  CMXI2X1 U24106 ( .A0(n13412), .A1(n13436), .S(n3276), .Z(N8581) );
  CMX2X1 U24107 ( .A0(N7963), .A1(N7962), .S(n3865), .Z(n13419) );
  CMX2X1 U24108 ( .A0(n13414), .A1(n13426), .S(n4307), .Z(n13442) );
  CMXI2X1 U24109 ( .A0(n13415), .A1(n13442), .S(n3273), .Z(N8582) );
  CMX2X1 U24110 ( .A0(N7962), .A1(N7961), .S(n3866), .Z(n13422) );
  CMX2X1 U24111 ( .A0(n13417), .A1(n13429), .S(n4307), .Z(n13445) );
  CMXI2X1 U24112 ( .A0(n13418), .A1(n13445), .S(n3273), .Z(N8583) );
  CMX2X1 U24113 ( .A0(N7961), .A1(N7960), .S(n3867), .Z(n13425) );
  CMXI2X1 U24114 ( .A0(n13425), .A1(n13419), .S(n4184), .Z(n13432) );
  CMX2X1 U24115 ( .A0(n13420), .A1(n13432), .S(n4307), .Z(n13448) );
  CMXI2X1 U24116 ( .A0(n13421), .A1(n13448), .S(n3273), .Z(N8584) );
  CMX2X1 U24117 ( .A0(N7960), .A1(N7959), .S(n3868), .Z(n13428) );
  CMXI2X1 U24118 ( .A0(n13428), .A1(n13422), .S(n4184), .Z(n13435) );
  CMX2X1 U24119 ( .A0(n13423), .A1(n13435), .S(n3790), .Z(n13451) );
  CMXI2X1 U24120 ( .A0(n13424), .A1(n13451), .S(n3273), .Z(N8585) );
  CMX2X1 U24121 ( .A0(N7959), .A1(N7958), .S(n3878), .Z(n13431) );
  CMXI2X1 U24122 ( .A0(n13431), .A1(n13425), .S(n4184), .Z(n13441) );
  CMX2X1 U24123 ( .A0(n13426), .A1(n13441), .S(n3810), .Z(n13454) );
  CMXI2X1 U24124 ( .A0(n13427), .A1(n13454), .S(n3273), .Z(N8586) );
  CMX2X1 U24125 ( .A0(N7958), .A1(N7957), .S(n3868), .Z(n13434) );
  CMXI2X1 U24126 ( .A0(n13434), .A1(n13428), .S(n4184), .Z(n13444) );
  CMX2X1 U24127 ( .A0(n13429), .A1(n13444), .S(n3811), .Z(n13457) );
  CMXI2X1 U24128 ( .A0(n13430), .A1(n13457), .S(n3273), .Z(N8587) );
  CMX2X1 U24129 ( .A0(N7957), .A1(N7956), .S(n3869), .Z(n13440) );
  CMXI2X1 U24130 ( .A0(n13440), .A1(n13431), .S(n4184), .Z(n13447) );
  CMX2X1 U24131 ( .A0(n13432), .A1(n13447), .S(n3812), .Z(n13460) );
  CMXI2X1 U24132 ( .A0(n13433), .A1(n13460), .S(n3274), .Z(N8588) );
  CMX2X1 U24133 ( .A0(N7956), .A1(N7955), .S(n3873), .Z(n13443) );
  CMXI2X1 U24134 ( .A0(n13443), .A1(n13434), .S(n4184), .Z(n13450) );
  CMX2X1 U24135 ( .A0(n13435), .A1(n13450), .S(n4306), .Z(n13463) );
  CMXI2X1 U24136 ( .A0(n13436), .A1(n13463), .S(n3347), .Z(N8589) );
  CMX2X1 U24137 ( .A0(N8235), .A1(N8234), .S(n3874), .Z(n13503) );
  CMXI2X1 U24138 ( .A0(n13503), .A1(n13437), .S(n4184), .Z(n13570) );
  CMX2X1 U24139 ( .A0(n13438), .A1(n13570), .S(n3771), .Z(n13703) );
  CMXI2X1 U24140 ( .A0(n13439), .A1(n13703), .S(n3340), .Z(N8310) );
  CMX2X1 U24141 ( .A0(N7955), .A1(N7954), .S(n3881), .Z(n13446) );
  CMXI2X1 U24142 ( .A0(n13446), .A1(n13440), .S(n4184), .Z(n13453) );
  CMX2X1 U24143 ( .A0(n13441), .A1(n13453), .S(n3812), .Z(n13466) );
  CMXI2X1 U24144 ( .A0(n13442), .A1(n13466), .S(n3433), .Z(N8590) );
  CMX2X1 U24145 ( .A0(N7954), .A1(N7953), .S(n3862), .Z(n13449) );
  CMXI2X1 U24146 ( .A0(n13449), .A1(n13443), .S(n4184), .Z(n13456) );
  CMX2X1 U24147 ( .A0(n13444), .A1(n13456), .S(n3772), .Z(n13469) );
  CMXI2X1 U24148 ( .A0(n13445), .A1(n13469), .S(n3432), .Z(N8591) );
  CMX2X1 U24149 ( .A0(N7953), .A1(N7952), .S(n3863), .Z(n13452) );
  CMXI2X1 U24150 ( .A0(n13452), .A1(n13446), .S(n4184), .Z(n13459) );
  CMX2X1 U24151 ( .A0(n13447), .A1(n13459), .S(n3773), .Z(n13475) );
  CMXI2X1 U24152 ( .A0(n13448), .A1(n13475), .S(n3430), .Z(N8592) );
  CMX2X1 U24153 ( .A0(N7952), .A1(N7951), .S(n3864), .Z(n13455) );
  CMXI2X1 U24154 ( .A0(n13455), .A1(n13449), .S(n4184), .Z(n13462) );
  CMX2X1 U24155 ( .A0(n13450), .A1(n13462), .S(n3774), .Z(n13478) );
  CMXI2X1 U24156 ( .A0(n13451), .A1(n13478), .S(n3428), .Z(N8593) );
  CMX2X1 U24157 ( .A0(N7951), .A1(N7950), .S(n3879), .Z(n13458) );
  CMXI2X1 U24158 ( .A0(n13458), .A1(n13452), .S(n4184), .Z(n13465) );
  CMX2X1 U24159 ( .A0(n13453), .A1(n13465), .S(n3775), .Z(n13481) );
  CMXI2X1 U24160 ( .A0(n13454), .A1(n13481), .S(n3429), .Z(N8594) );
  CMX2X1 U24161 ( .A0(N7950), .A1(N7949), .S(n3880), .Z(n13461) );
  CMXI2X1 U24162 ( .A0(n13461), .A1(n13455), .S(n4183), .Z(n13468) );
  CMX2X1 U24163 ( .A0(n13456), .A1(n13468), .S(n4306), .Z(n13484) );
  CMXI2X1 U24164 ( .A0(n13457), .A1(n13484), .S(n3333), .Z(N8595) );
  CMX2X1 U24165 ( .A0(N7949), .A1(N7948), .S(n3881), .Z(n13464) );
  CMXI2X1 U24166 ( .A0(n13464), .A1(n13458), .S(n4183), .Z(n13474) );
  CMX2X1 U24167 ( .A0(n13459), .A1(n13474), .S(n4306), .Z(n13487) );
  CMXI2X1 U24168 ( .A0(n13460), .A1(n13487), .S(n3333), .Z(N8596) );
  CMX2X1 U24169 ( .A0(N7948), .A1(N7947), .S(n3862), .Z(n13467) );
  CMXI2X1 U24170 ( .A0(n13467), .A1(n13461), .S(n4183), .Z(n13477) );
  CMX2X1 U24171 ( .A0(n13462), .A1(n13477), .S(n4306), .Z(n13490) );
  CMXI2X1 U24172 ( .A0(n13463), .A1(n13490), .S(n3333), .Z(N8597) );
  CMX2X1 U24173 ( .A0(N7947), .A1(N7946), .S(n3871), .Z(n13473) );
  CMXI2X1 U24174 ( .A0(n13473), .A1(n13464), .S(n4183), .Z(n13480) );
  CMX2X1 U24175 ( .A0(n13465), .A1(n13480), .S(n4306), .Z(n13493) );
  CMXI2X1 U24176 ( .A0(n13466), .A1(n13493), .S(n3333), .Z(N8598) );
  CMX2X1 U24177 ( .A0(N7946), .A1(N7945), .S(n3875), .Z(n13476) );
  CMXI2X1 U24178 ( .A0(n13476), .A1(n13467), .S(n4183), .Z(n13483) );
  CMX2X1 U24179 ( .A0(n13468), .A1(n13483), .S(n4306), .Z(n13496) );
  CMXI2X1 U24180 ( .A0(n13469), .A1(n13496), .S(n3333), .Z(N8599) );
  CMX2X1 U24181 ( .A0(N8234), .A1(N8233), .S(n3876), .Z(n13536) );
  CMXI2X1 U24182 ( .A0(n13536), .A1(n13470), .S(n4183), .Z(n13603) );
  CMX2X1 U24183 ( .A0(n13471), .A1(n13603), .S(n4306), .Z(n13736) );
  CMXI2X1 U24184 ( .A0(n13472), .A1(n13736), .S(n3333), .Z(N8311) );
  CMX2X1 U24185 ( .A0(N7945), .A1(N7944), .S(n3877), .Z(n13479) );
  CMXI2X1 U24186 ( .A0(n13479), .A1(n13473), .S(n4183), .Z(n13486) );
  CMX2X1 U24187 ( .A0(n13474), .A1(n13486), .S(n4306), .Z(n13499) );
  CMXI2X1 U24188 ( .A0(n13475), .A1(n13499), .S(n3333), .Z(N8600) );
  CMX2X1 U24189 ( .A0(N7944), .A1(N7943), .S(n3878), .Z(n13482) );
  CMXI2X1 U24190 ( .A0(n13482), .A1(n13476), .S(n4183), .Z(n13489) );
  CMX2X1 U24191 ( .A0(n13477), .A1(n13489), .S(n4306), .Z(n13502) );
  CMXI2X1 U24192 ( .A0(n13478), .A1(n13502), .S(n3335), .Z(N8601) );
  CMX2X1 U24193 ( .A0(N7943), .A1(N7942), .S(n3879), .Z(n13485) );
  CMXI2X1 U24194 ( .A0(n13485), .A1(n13479), .S(n4183), .Z(n13492) );
  CMX2X1 U24195 ( .A0(n13480), .A1(n13492), .S(n4306), .Z(n13508) );
  CMXI2X1 U24196 ( .A0(n13481), .A1(n13508), .S(n3335), .Z(N8602) );
  CMX2X1 U24197 ( .A0(N7942), .A1(N7941), .S(n3880), .Z(n13488) );
  CMX2X1 U24198 ( .A0(n13483), .A1(n13495), .S(n4306), .Z(n13511) );
  CMXI2X1 U24199 ( .A0(n13484), .A1(n13511), .S(n3335), .Z(N8603) );
  CMX2X1 U24200 ( .A0(N7941), .A1(N7940), .S(n3881), .Z(n13491) );
  CMXI2X1 U24201 ( .A0(n13491), .A1(n13485), .S(n4183), .Z(n13498) );
  CMX2X1 U24202 ( .A0(n13486), .A1(n13498), .S(n4306), .Z(n13514) );
  CMXI2X1 U24203 ( .A0(n13487), .A1(n13514), .S(n3335), .Z(N8604) );
  CMX2X1 U24204 ( .A0(N7940), .A1(N7939), .S(n3870), .Z(n13494) );
  CMXI2X1 U24205 ( .A0(n13494), .A1(n13488), .S(n4183), .Z(n13501) );
  CMX2X1 U24206 ( .A0(n13489), .A1(n13501), .S(n4305), .Z(n13517) );
  CMXI2X1 U24207 ( .A0(n13490), .A1(n13517), .S(n3335), .Z(N8605) );
  CMX2X1 U24208 ( .A0(N7939), .A1(N7938), .S(n3871), .Z(n13497) );
  CMXI2X1 U24209 ( .A0(n13497), .A1(n13491), .S(n4183), .Z(n13507) );
  CMX2X1 U24210 ( .A0(n13492), .A1(n13507), .S(n4305), .Z(n13520) );
  CMXI2X1 U24211 ( .A0(n13493), .A1(n13520), .S(n3335), .Z(N8606) );
  CMX2X1 U24212 ( .A0(N7938), .A1(N7937), .S(n3862), .Z(n13500) );
  CMXI2X1 U24213 ( .A0(n13500), .A1(n13494), .S(n4183), .Z(n13510) );
  CMX2X1 U24214 ( .A0(n13495), .A1(n13510), .S(n4305), .Z(n13523) );
  CMXI2X1 U24215 ( .A0(n13496), .A1(n13523), .S(n3335), .Z(N8607) );
  CMX2X1 U24216 ( .A0(N7937), .A1(N7936), .S(n3863), .Z(n13506) );
  CMXI2X1 U24217 ( .A0(n13506), .A1(n13497), .S(n4183), .Z(n13513) );
  CMX2X1 U24218 ( .A0(n13498), .A1(n13513), .S(n4305), .Z(n13526) );
  CMXI2X1 U24219 ( .A0(n13499), .A1(n13526), .S(n3334), .Z(N8608) );
  CMX2X1 U24220 ( .A0(N7936), .A1(N7935), .S(n3865), .Z(n13509) );
  CMXI2X1 U24221 ( .A0(n13509), .A1(n13500), .S(n4183), .Z(n13516) );
  CMX2X1 U24222 ( .A0(n13501), .A1(n13516), .S(n4305), .Z(n13529) );
  CMXI2X1 U24223 ( .A0(n13502), .A1(n13529), .S(n3334), .Z(N8609) );
  CMX2X1 U24224 ( .A0(N8233), .A1(N8232), .S(n3866), .Z(n13569) );
  CMXI2X1 U24225 ( .A0(n13569), .A1(n13503), .S(n4182), .Z(n13636) );
  CMX2X1 U24226 ( .A0(n13504), .A1(n13636), .S(n4305), .Z(n13776) );
  CMXI2X1 U24227 ( .A0(n13505), .A1(n13776), .S(n3334), .Z(N8312) );
  CMX2X1 U24228 ( .A0(N7935), .A1(N7934), .S(n3867), .Z(n13512) );
  CMXI2X1 U24229 ( .A0(n13512), .A1(n13506), .S(n4182), .Z(n13519) );
  CMX2X1 U24230 ( .A0(n13507), .A1(n13519), .S(n4305), .Z(n13532) );
  CMXI2X1 U24231 ( .A0(n13508), .A1(n13532), .S(n3334), .Z(N8610) );
  CMX2X1 U24232 ( .A0(N7934), .A1(N7933), .S(n3868), .Z(n13515) );
  CMXI2X1 U24233 ( .A0(n13515), .A1(n13509), .S(n4182), .Z(n13522) );
  CMX2X1 U24234 ( .A0(n13510), .A1(n13522), .S(n4305), .Z(n13535) );
  CMXI2X1 U24235 ( .A0(n13511), .A1(n13535), .S(n3334), .Z(N8611) );
  CMX2X1 U24236 ( .A0(N7933), .A1(N7932), .S(n3863), .Z(n13518) );
  CMXI2X1 U24237 ( .A0(n13518), .A1(n13512), .S(n4182), .Z(n13525) );
  CMX2X1 U24238 ( .A0(n13513), .A1(n13525), .S(n4305), .Z(n13541) );
  CMXI2X1 U24239 ( .A0(n13514), .A1(n13541), .S(n3334), .Z(N8612) );
  CMX2X1 U24240 ( .A0(N7932), .A1(N7931), .S(n3864), .Z(n13521) );
  CMXI2X1 U24241 ( .A0(n13521), .A1(n13515), .S(n4182), .Z(n13528) );
  CMX2X1 U24242 ( .A0(n13516), .A1(n13528), .S(n4305), .Z(n13544) );
  CMXI2X1 U24243 ( .A0(n13517), .A1(n13544), .S(n3334), .Z(N8613) );
  CMX2X1 U24244 ( .A0(N7931), .A1(N7930), .S(n3865), .Z(n13524) );
  CMXI2X1 U24245 ( .A0(n13524), .A1(n13518), .S(n4182), .Z(n13531) );
  CMX2X1 U24246 ( .A0(n13519), .A1(n13531), .S(n4305), .Z(n13547) );
  CMXI2X1 U24247 ( .A0(n13520), .A1(n13547), .S(n3334), .Z(N8614) );
  CMX2X1 U24248 ( .A0(N7930), .A1(N7929), .S(n3866), .Z(n13527) );
  CMX2X1 U24249 ( .A0(n13522), .A1(n13534), .S(n3812), .Z(n13550) );
  CMXI2X1 U24250 ( .A0(n13523), .A1(n13550), .S(n3334), .Z(N8615) );
  CMX2X1 U24251 ( .A0(N7929), .A1(N7928), .S(n3872), .Z(n13530) );
  CMXI2X1 U24252 ( .A0(n13530), .A1(n13524), .S(n4182), .Z(n13540) );
  CMX2X1 U24253 ( .A0(n13525), .A1(n13540), .S(n4375), .Z(n13553) );
  CMXI2X1 U24254 ( .A0(n13526), .A1(n13553), .S(n3334), .Z(N8616) );
  CMX2X1 U24255 ( .A0(N7928), .A1(N7927), .S(n3864), .Z(n13533) );
  CMXI2X1 U24256 ( .A0(n13533), .A1(n13527), .S(n4182), .Z(n13543) );
  CMX2X1 U24257 ( .A0(n13528), .A1(n13543), .S(n3794), .Z(n13556) );
  CMXI2X1 U24258 ( .A0(n13529), .A1(n13556), .S(n3334), .Z(N8617) );
  CMX2X1 U24259 ( .A0(N7927), .A1(N7926), .S(n3865), .Z(n13539) );
  CMXI2X1 U24260 ( .A0(n13539), .A1(n13530), .S(n4182), .Z(n13546) );
  CMX2X1 U24261 ( .A0(n13531), .A1(n13546), .S(n3795), .Z(n13559) );
  CMXI2X1 U24262 ( .A0(n13532), .A1(n13559), .S(n3337), .Z(N8618) );
  CMX2X1 U24263 ( .A0(N7926), .A1(N7925), .S(n3866), .Z(n13542) );
  CMX2X1 U24264 ( .A0(n13534), .A1(n13549), .S(n3796), .Z(n13562) );
  CMXI2X1 U24265 ( .A0(n13535), .A1(n13562), .S(n3337), .Z(N8619) );
  CMX2X1 U24266 ( .A0(N8232), .A1(N8231), .S(n3867), .Z(n13602) );
  CMXI2X1 U24267 ( .A0(n13602), .A1(n13536), .S(n4182), .Z(n13669) );
  CMX2X1 U24268 ( .A0(n13537), .A1(n13669), .S(n3797), .Z(n13809) );
  CMXI2X1 U24269 ( .A0(n13538), .A1(n13809), .S(n3336), .Z(N8313) );
  CMX2X1 U24270 ( .A0(N7925), .A1(N7924), .S(n3868), .Z(n13545) );
  CMX2X1 U24271 ( .A0(n13540), .A1(n13552), .S(n3805), .Z(n13565) );
  CMXI2X1 U24272 ( .A0(n13541), .A1(n13565), .S(n3336), .Z(N8620) );
  CMX2X1 U24273 ( .A0(N7924), .A1(N7923), .S(n3869), .Z(n13548) );
  CMXI2X1 U24274 ( .A0(n13548), .A1(n13542), .S(n4182), .Z(n13555) );
  CMX2X1 U24275 ( .A0(n13543), .A1(n13555), .S(n3809), .Z(n13568) );
  CMXI2X1 U24276 ( .A0(n13544), .A1(n13568), .S(n3336), .Z(N8621) );
  CMX2X1 U24277 ( .A0(N7923), .A1(N7922), .S(n3870), .Z(n13551) );
  CMXI2X1 U24278 ( .A0(n13551), .A1(n13545), .S(n4182), .Z(n13558) );
  CMX2X1 U24279 ( .A0(n13546), .A1(n13558), .S(n3772), .Z(n13574) );
  CMXI2X1 U24280 ( .A0(n13547), .A1(n13574), .S(n3336), .Z(N8622) );
  CMX2X1 U24281 ( .A0(N7922), .A1(N7921), .S(n3872), .Z(n13554) );
  CMXI2X1 U24282 ( .A0(n13554), .A1(n13548), .S(n4182), .Z(n13561) );
  CMX2X1 U24283 ( .A0(n13549), .A1(n13561), .S(n3773), .Z(n13577) );
  CMXI2X1 U24284 ( .A0(n13550), .A1(n13577), .S(n3336), .Z(N8623) );
  CMX2X1 U24285 ( .A0(N7921), .A1(N7920), .S(n3873), .Z(n13557) );
  CMXI2X1 U24286 ( .A0(n13557), .A1(n13551), .S(n4181), .Z(n13564) );
  CMX2X1 U24287 ( .A0(n13552), .A1(n13564), .S(n3774), .Z(n13580) );
  CMXI2X1 U24288 ( .A0(n13553), .A1(n13580), .S(n3336), .Z(N8624) );
  CMX2X1 U24289 ( .A0(N7920), .A1(N7919), .S(n3871), .Z(n13560) );
  CMXI2X1 U24290 ( .A0(n13560), .A1(n13554), .S(n4181), .Z(n13567) );
  CMX2X1 U24291 ( .A0(n13555), .A1(n13567), .S(n3797), .Z(n13583) );
  CMXI2X1 U24292 ( .A0(n13556), .A1(n13583), .S(n3336), .Z(N8625) );
  CMX2X1 U24293 ( .A0(N7919), .A1(N7918), .S(n3872), .Z(n13563) );
  CMXI2X1 U24294 ( .A0(n13563), .A1(n13557), .S(n4181), .Z(n13573) );
  CMX2X1 U24295 ( .A0(n13558), .A1(n13573), .S(n3805), .Z(n13586) );
  CMXI2X1 U24296 ( .A0(n13559), .A1(n13586), .S(n3336), .Z(N8626) );
  CMX2X1 U24297 ( .A0(N7918), .A1(N7917), .S(n3869), .Z(n13566) );
  CMXI2X1 U24298 ( .A0(n13566), .A1(n13560), .S(n4181), .Z(n13576) );
  CMX2X1 U24299 ( .A0(n13561), .A1(n13576), .S(n3806), .Z(n13589) );
  CMXI2X1 U24300 ( .A0(n13562), .A1(n13589), .S(n3336), .Z(N8627) );
  CMX2X1 U24301 ( .A0(N7917), .A1(N7916), .S(n3870), .Z(n13572) );
  CMX2X1 U24302 ( .A0(n13564), .A1(n3709), .S(n3807), .Z(n13592) );
  CMXI2X1 U24303 ( .A0(n13565), .A1(n13592), .S(n3336), .Z(N8628) );
  CMX2X1 U24304 ( .A0(N7916), .A1(N7915), .S(n3871), .Z(n13575) );
  CMXI2X1 U24305 ( .A0(n13575), .A1(n13566), .S(n4181), .Z(n13582) );
  CMX2X1 U24306 ( .A0(n13567), .A1(n13582), .S(n3808), .Z(n13595) );
  CMXI2X1 U24307 ( .A0(n13568), .A1(n13595), .S(n3336), .Z(N8629) );
  CMX2X1 U24308 ( .A0(N8231), .A1(N8230), .S(n3872), .Z(n13635) );
  CMXI2X1 U24309 ( .A0(n13635), .A1(n13569), .S(n4181), .Z(n13702) );
  CMX2X1 U24310 ( .A0(n13570), .A1(n13702), .S(n3809), .Z(n13842) );
  CMXI2X1 U24311 ( .A0(n13571), .A1(n13842), .S(n3335), .Z(N8314) );
  CMX2X1 U24312 ( .A0(N7915), .A1(N7914), .S(n3867), .Z(n13578) );
  CMXI2X1 U24313 ( .A0(n13578), .A1(n13572), .S(n4181), .Z(n13585) );
  CMX2X1 U24314 ( .A0(n13573), .A1(n13585), .S(n3810), .Z(n13598) );
  CMXI2X1 U24315 ( .A0(n13574), .A1(n13598), .S(n3335), .Z(N8630) );
  CMX2X1 U24316 ( .A0(N7914), .A1(N7913), .S(n3868), .Z(n13581) );
  CMXI2X1 U24317 ( .A0(n13581), .A1(n13575), .S(n4181), .Z(n13588) );
  CMX2X1 U24318 ( .A0(n13576), .A1(n13588), .S(n3811), .Z(n13601) );
  CMXI2X1 U24319 ( .A0(n13577), .A1(n13601), .S(n3335), .Z(N8631) );
  CMX2X1 U24320 ( .A0(N7913), .A1(N7912), .S(n3869), .Z(n13584) );
  CMXI2X1 U24321 ( .A0(n13584), .A1(n13578), .S(n4181), .Z(n13591) );
  CMX2X1 U24322 ( .A0(n13579), .A1(n13591), .S(n3812), .Z(n13607) );
  CMXI2X1 U24323 ( .A0(n13580), .A1(n13607), .S(n3335), .Z(N8632) );
  CMX2X1 U24324 ( .A0(N7912), .A1(N7911), .S(n3870), .Z(n13587) );
  CMXI2X1 U24325 ( .A0(n13587), .A1(n13581), .S(n4181), .Z(n13594) );
  CMX2X1 U24326 ( .A0(n13582), .A1(n13594), .S(n4305), .Z(n13610) );
  CMX2X1 U24327 ( .A0(N7911), .A1(N7910), .S(n3873), .Z(n13590) );
  CMXI2X1 U24328 ( .A0(n13590), .A1(n13584), .S(n4181), .Z(n13597) );
  CMX2X1 U24329 ( .A0(n13585), .A1(n13597), .S(n3771), .Z(n13613) );
  CMX2X1 U24330 ( .A0(N7910), .A1(N7909), .S(n3873), .Z(n13593) );
  CMXI2X1 U24331 ( .A0(n13593), .A1(n13587), .S(n4181), .Z(n13600) );
  CMX2X1 U24332 ( .A0(n13588), .A1(n13600), .S(n3777), .Z(n13616) );
  CMXI2X1 U24333 ( .A0(n13589), .A1(n13616), .S(n3338), .Z(N8635) );
  CMX2X1 U24334 ( .A0(N7909), .A1(N7908), .S(n3874), .Z(n13596) );
  CMXI2X1 U24335 ( .A0(n13596), .A1(n13590), .S(n4181), .Z(n13606) );
  CMX2X1 U24336 ( .A0(n13591), .A1(n13606), .S(n3790), .Z(n13619) );
  CMXI2X1 U24337 ( .A0(n13592), .A1(n13619), .S(n3338), .Z(N8636) );
  CMX2X1 U24338 ( .A0(N7908), .A1(N7907), .S(n3875), .Z(n13599) );
  CMXI2X1 U24339 ( .A0(n13599), .A1(n13593), .S(n4181), .Z(n13609) );
  CMX2X1 U24340 ( .A0(n13594), .A1(n13609), .S(n3791), .Z(n13622) );
  CMXI2X1 U24341 ( .A0(n13595), .A1(n13622), .S(n3338), .Z(N8637) );
  CMX2X1 U24342 ( .A0(N7907), .A1(N7906), .S(n3876), .Z(n13605) );
  CMXI2X1 U24343 ( .A0(n13605), .A1(n13596), .S(n4181), .Z(n13612) );
  CMX2X1 U24344 ( .A0(n13597), .A1(n13612), .S(n3792), .Z(n13625) );
  CMXI2X1 U24345 ( .A0(n13598), .A1(n13625), .S(n3338), .Z(N8638) );
  CMX2X1 U24346 ( .A0(N7906), .A1(N7905), .S(n3877), .Z(n13608) );
  CMXI2X1 U24347 ( .A0(n13608), .A1(n13599), .S(n4180), .Z(n13615) );
  CMX2X1 U24348 ( .A0(n13600), .A1(n13615), .S(n3793), .Z(n13628) );
  CMX2X1 U24349 ( .A0(N8230), .A1(N8229), .S(n3878), .Z(n13668) );
  CMXI2X1 U24350 ( .A0(n13668), .A1(n13602), .S(n4180), .Z(n13735) );
  CMX2X1 U24351 ( .A0(n13603), .A1(n13735), .S(n3808), .Z(n13874) );
  CMXI2X1 U24352 ( .A0(n13604), .A1(n13874), .S(n3338), .Z(N8315) );
  CMX2X1 U24353 ( .A0(N7905), .A1(N7904), .S(n3879), .Z(n13611) );
  CMXI2X1 U24354 ( .A0(n13611), .A1(n13605), .S(n4180), .Z(n13618) );
  CMX2X1 U24355 ( .A0(n13606), .A1(n13618), .S(n3792), .Z(n13631) );
  CMXI2X1 U24356 ( .A0(n13607), .A1(n13631), .S(n3338), .Z(N8640) );
  CMX2X1 U24357 ( .A0(N7904), .A1(N7903), .S(n3874), .Z(n13614) );
  CMXI2X1 U24358 ( .A0(n13614), .A1(n13608), .S(n4180), .Z(n13621) );
  CMX2X1 U24359 ( .A0(n13609), .A1(n13621), .S(n3793), .Z(n13634) );
  CMXI2X1 U24360 ( .A0(n13610), .A1(n13634), .S(n3338), .Z(N8641) );
  CMX2X1 U24361 ( .A0(N7903), .A1(N7902), .S(n3875), .Z(n13617) );
  CMXI2X1 U24362 ( .A0(n13617), .A1(n13611), .S(n4180), .Z(n13624) );
  CMX2X1 U24363 ( .A0(n13612), .A1(n13624), .S(n3794), .Z(n13640) );
  CMXI2X1 U24364 ( .A0(n13613), .A1(n13640), .S(n3337), .Z(N8642) );
  CMX2X1 U24365 ( .A0(N7902), .A1(N7901), .S(n3880), .Z(n13620) );
  CMX2X1 U24366 ( .A0(n13615), .A1(n13627), .S(n3795), .Z(n13643) );
  CMXI2X1 U24367 ( .A0(n13616), .A1(n13643), .S(n3337), .Z(N8643) );
  CMX2X1 U24368 ( .A0(N7901), .A1(N7900), .S(n3881), .Z(n13623) );
  CMXI2X1 U24369 ( .A0(n13623), .A1(n13617), .S(n4180), .Z(n13630) );
  CMX2X1 U24370 ( .A0(n13618), .A1(n13630), .S(n3796), .Z(n13646) );
  CMXI2X1 U24371 ( .A0(n13619), .A1(n13646), .S(n3337), .Z(N8644) );
  CMX2X1 U24372 ( .A0(N7900), .A1(N7899), .S(n3873), .Z(n13626) );
  CMXI2X1 U24373 ( .A0(n13626), .A1(n13620), .S(n4180), .Z(n13633) );
  CMX2X1 U24374 ( .A0(n13621), .A1(n13633), .S(n3771), .Z(n13649) );
  CMXI2X1 U24375 ( .A0(n13622), .A1(n13649), .S(n3337), .Z(N8645) );
  CMX2X1 U24376 ( .A0(N7899), .A1(N7898), .S(n3874), .Z(n13629) );
  CMXI2X1 U24377 ( .A0(n13629), .A1(n13623), .S(n4180), .Z(n13639) );
  CMX2X1 U24378 ( .A0(n13624), .A1(n13639), .S(n3772), .Z(n13652) );
  CMXI2X1 U24379 ( .A0(n13625), .A1(n13652), .S(n3337), .Z(N8646) );
  CMX2X1 U24380 ( .A0(N7898), .A1(N7897), .S(n3875), .Z(n13632) );
  CMXI2X1 U24381 ( .A0(n13632), .A1(n13626), .S(n4180), .Z(n13642) );
  CMX2X1 U24382 ( .A0(n13627), .A1(n13642), .S(n3773), .Z(n13655) );
  CMXI2X1 U24383 ( .A0(n13628), .A1(n13655), .S(n3337), .Z(N8647) );
  CMX2X1 U24384 ( .A0(N7897), .A1(N7896), .S(n3876), .Z(n13638) );
  CMXI2X1 U24385 ( .A0(n13638), .A1(n13629), .S(n4180), .Z(n13645) );
  CMX2X1 U24386 ( .A0(n3708), .A1(n13645), .S(n3774), .Z(n13658) );
  CMXI2X1 U24387 ( .A0(n13631), .A1(n13658), .S(n3337), .Z(N8648) );
  CMX2X1 U24388 ( .A0(N7896), .A1(N7895), .S(n3872), .Z(n13641) );
  CMXI2X1 U24389 ( .A0(n13641), .A1(n13632), .S(n4180), .Z(n13648) );
  CMX2X1 U24390 ( .A0(n13633), .A1(n13648), .S(n3775), .Z(n13661) );
  CMXI2X1 U24391 ( .A0(n13634), .A1(n13661), .S(n3337), .Z(N8649) );
  CMX2X1 U24392 ( .A0(N8229), .A1(N8228), .S(n3873), .Z(n13701) );
  CMXI2X1 U24393 ( .A0(n13701), .A1(n13635), .S(n4180), .Z(n13775) );
  CMX2X1 U24394 ( .A0(n13636), .A1(n13775), .S(n3776), .Z(n13907) );
  CMXI2X1 U24395 ( .A0(n13637), .A1(n13907), .S(n3337), .Z(N8316) );
  CMX2X1 U24396 ( .A0(N7895), .A1(N7894), .S(n3874), .Z(n13644) );
  CMXI2X1 U24397 ( .A0(n13644), .A1(n13638), .S(n4180), .Z(n13651) );
  CMX2X1 U24398 ( .A0(n13639), .A1(n13651), .S(n3777), .Z(n13664) );
  CMXI2X1 U24399 ( .A0(n13640), .A1(n13664), .S(n3340), .Z(N8650) );
  CMX2X1 U24400 ( .A0(N7894), .A1(N7893), .S(n3874), .Z(n13647) );
  CMXI2X1 U24401 ( .A0(n13647), .A1(n13641), .S(n4180), .Z(n13654) );
  CMX2X1 U24402 ( .A0(n13642), .A1(n13654), .S(n3790), .Z(n13667) );
  CMXI2X1 U24403 ( .A0(n13643), .A1(n13667), .S(n3339), .Z(N8651) );
  CMX2X1 U24404 ( .A0(N7893), .A1(N7892), .S(n3862), .Z(n13650) );
  CMXI2X1 U24405 ( .A0(n13650), .A1(n13644), .S(n4180), .Z(n13657) );
  CMX2X1 U24406 ( .A0(n13645), .A1(n13657), .S(n3791), .Z(n13673) );
  CMXI2X1 U24407 ( .A0(n13646), .A1(n13673), .S(n3339), .Z(N8652) );
  CMX2X1 U24408 ( .A0(N7892), .A1(N7891), .S(n3863), .Z(n13653) );
  CMXI2X1 U24409 ( .A0(n13653), .A1(n13647), .S(n4179), .Z(n13660) );
  CMX2X1 U24410 ( .A0(n13648), .A1(n13660), .S(n3811), .Z(n13676) );
  CMXI2X1 U24411 ( .A0(n13649), .A1(n13676), .S(n3339), .Z(N8653) );
  CMX2X1 U24412 ( .A0(N7891), .A1(N7890), .S(n3864), .Z(n13656) );
  CMXI2X1 U24413 ( .A0(n13656), .A1(n13650), .S(n4179), .Z(n13663) );
  CMX2X1 U24414 ( .A0(n13651), .A1(n13663), .S(n3812), .Z(n13679) );
  CMX2X1 U24415 ( .A0(N7890), .A1(N7889), .S(n3865), .Z(n13659) );
  CMX2X1 U24416 ( .A0(n13654), .A1(n13666), .S(n3774), .Z(n13682) );
  CMXI2X1 U24417 ( .A0(n13655), .A1(n13682), .S(n3339), .Z(N8655) );
  CMX2X1 U24418 ( .A0(N7889), .A1(N7888), .S(n3866), .Z(n13662) );
  CMXI2X1 U24419 ( .A0(n13662), .A1(n13656), .S(n4179), .Z(n13672) );
  CMX2X1 U24420 ( .A0(n13657), .A1(n13672), .S(n3775), .Z(n13685) );
  CMXI2X1 U24421 ( .A0(n13658), .A1(n13685), .S(n3339), .Z(N8656) );
  CMX2X1 U24422 ( .A0(N7888), .A1(N7887), .S(n3867), .Z(n13665) );
  CMXI2X1 U24423 ( .A0(n13665), .A1(n13659), .S(n4179), .Z(n13675) );
  CMX2X1 U24424 ( .A0(n13660), .A1(n13675), .S(n3776), .Z(n13688) );
  CMXI2X1 U24425 ( .A0(n13661), .A1(n13688), .S(n3339), .Z(N8657) );
  CMX2X1 U24426 ( .A0(N7887), .A1(N7886), .S(n3868), .Z(n13671) );
  CMXI2X1 U24427 ( .A0(n13671), .A1(n13662), .S(n4179), .Z(n13678) );
  CMX2X1 U24428 ( .A0(n13663), .A1(n13678), .S(n3807), .Z(n13691) );
  CMX2X1 U24429 ( .A0(N7886), .A1(N7885), .S(n3876), .Z(n13674) );
  CMXI2X1 U24430 ( .A0(n13674), .A1(n13665), .S(n4179), .Z(n13681) );
  CMX2X1 U24431 ( .A0(n13666), .A1(n13681), .S(n3807), .Z(n13694) );
  CMXI2X1 U24432 ( .A0(n13667), .A1(n13694), .S(n3339), .Z(N8659) );
  CMX2X1 U24433 ( .A0(N8228), .A1(N8227), .S(n3877), .Z(n13734) );
  CMXI2X1 U24434 ( .A0(n13734), .A1(n13668), .S(n4179), .Z(n13808) );
  CMX2X1 U24435 ( .A0(n13669), .A1(n13808), .S(n3808), .Z(n13940) );
  CMXI2X1 U24436 ( .A0(n13670), .A1(n13940), .S(n3339), .Z(N8317) );
  CMX2X1 U24437 ( .A0(N7885), .A1(N7884), .S(n3869), .Z(n13677) );
  CMXI2X1 U24438 ( .A0(n13677), .A1(n13671), .S(n4179), .Z(n13684) );
  CMX2X1 U24439 ( .A0(n13672), .A1(n13684), .S(n3809), .Z(n13697) );
  CMXI2X1 U24440 ( .A0(n13673), .A1(n13697), .S(n3339), .Z(N8660) );
  CMX2X1 U24441 ( .A0(N7884), .A1(N7883), .S(n3870), .Z(n13680) );
  CMXI2X1 U24442 ( .A0(n13680), .A1(n13674), .S(n4179), .Z(n13687) );
  CMX2X1 U24443 ( .A0(n13675), .A1(n13687), .S(n3810), .Z(n13700) );
  CMXI2X1 U24444 ( .A0(n13676), .A1(n13700), .S(n3339), .Z(N8661) );
  CMX2X1 U24445 ( .A0(N7883), .A1(N7882), .S(n3877), .Z(n13683) );
  CMXI2X1 U24446 ( .A0(n13683), .A1(n13677), .S(n4179), .Z(n13690) );
  CMX2X1 U24447 ( .A0(n13678), .A1(n13690), .S(n3812), .Z(n13706) );
  CMXI2X1 U24448 ( .A0(n13679), .A1(n13706), .S(n3339), .Z(N8662) );
  CMX2X1 U24449 ( .A0(N7882), .A1(N7881), .S(n3878), .Z(n13686) );
  CMXI2X1 U24450 ( .A0(n13686), .A1(n13680), .S(n4179), .Z(n13693) );
  CMX2X1 U24451 ( .A0(n13681), .A1(n13693), .S(n4372), .Z(n13709) );
  CMXI2X1 U24452 ( .A0(n13682), .A1(n13709), .S(n3338), .Z(N8663) );
  CMX2X1 U24453 ( .A0(N7881), .A1(N7880), .S(n3879), .Z(n13689) );
  CMXI2X1 U24454 ( .A0(n13689), .A1(n13683), .S(n4179), .Z(n13696) );
  CMX2X1 U24455 ( .A0(n13684), .A1(n13696), .S(n3793), .Z(n13712) );
  CMXI2X1 U24456 ( .A0(n13685), .A1(n13712), .S(n3338), .Z(N8664) );
  CMX2X1 U24457 ( .A0(N7880), .A1(N7879), .S(n3880), .Z(n13692) );
  CMXI2X1 U24458 ( .A0(n13692), .A1(n13686), .S(n4179), .Z(n13699) );
  CMX2X1 U24459 ( .A0(n13687), .A1(n13699), .S(n3794), .Z(n13715) );
  CMXI2X1 U24460 ( .A0(n13688), .A1(n13715), .S(n3338), .Z(N8665) );
  CMX2X1 U24461 ( .A0(N7879), .A1(N7878), .S(n3875), .Z(n13695) );
  CMXI2X1 U24462 ( .A0(n13695), .A1(n13689), .S(n4179), .Z(n13705) );
  CMX2X1 U24463 ( .A0(n13690), .A1(n13705), .S(n3795), .Z(n13718) );
  CMXI2X1 U24464 ( .A0(n13691), .A1(n13718), .S(n3338), .Z(N8666) );
  CMX2X1 U24465 ( .A0(N7878), .A1(N7877), .S(n3876), .Z(n13698) );
  CMXI2X1 U24466 ( .A0(n13698), .A1(n13692), .S(n4179), .Z(n13708) );
  CMX2X1 U24467 ( .A0(n13693), .A1(n13708), .S(n3796), .Z(n13721) );
  CMXI2X1 U24468 ( .A0(n13694), .A1(n13721), .S(n3341), .Z(N8667) );
  CMX2X1 U24469 ( .A0(N7877), .A1(N7876), .S(n3877), .Z(n13704) );
  CMXI2X1 U24470 ( .A0(n13704), .A1(n13695), .S(n4178), .Z(n13711) );
  CMX2X1 U24471 ( .A0(n13696), .A1(n13711), .S(n3797), .Z(n13724) );
  CMXI2X1 U24472 ( .A0(n13697), .A1(n13724), .S(n3341), .Z(N8668) );
  CMX2X1 U24473 ( .A0(N7876), .A1(N7875), .S(n3878), .Z(n13707) );
  CMXI2X1 U24474 ( .A0(n13707), .A1(n13698), .S(n4178), .Z(n13714) );
  CMX2X1 U24475 ( .A0(n13699), .A1(n13714), .S(n3805), .Z(n13727) );
  CMXI2X1 U24476 ( .A0(n13700), .A1(n13727), .S(n3341), .Z(N8669) );
  CMX2X1 U24477 ( .A0(N8227), .A1(N8226), .S(n3875), .Z(n13774) );
  CMXI2X1 U24478 ( .A0(n13774), .A1(n13701), .S(n4178), .Z(n13841) );
  CMX2X1 U24479 ( .A0(n13702), .A1(n13841), .S(n3806), .Z(n13973) );
  CMXI2X1 U24480 ( .A0(n13703), .A1(n13973), .S(n3341), .Z(N8318) );
  CMX2X1 U24481 ( .A0(N7875), .A1(N7874), .S(n3871), .Z(n13710) );
  CMXI2X1 U24482 ( .A0(n13710), .A1(n13704), .S(n4178), .Z(n13717) );
  CMX2X1 U24483 ( .A0(n13705), .A1(n13717), .S(n3810), .Z(n13730) );
  CMXI2X1 U24484 ( .A0(n13706), .A1(n13730), .S(n3341), .Z(N8670) );
  CMX2X1 U24485 ( .A0(N7874), .A1(N7873), .S(n3872), .Z(n13713) );
  CMXI2X1 U24486 ( .A0(n13713), .A1(n13707), .S(n4178), .Z(n13720) );
  CMX2X1 U24487 ( .A0(n13708), .A1(n13720), .S(n3811), .Z(n13733) );
  CMXI2X1 U24488 ( .A0(n13709), .A1(n13733), .S(n3341), .Z(N8671) );
  CMX2X1 U24489 ( .A0(N7873), .A1(N7872), .S(n3873), .Z(n13716) );
  CMXI2X1 U24490 ( .A0(n13716), .A1(n13710), .S(n4178), .Z(n13723) );
  CMX2X1 U24491 ( .A0(n13711), .A1(n13723), .S(n3772), .Z(n13746) );
  CMXI2X1 U24492 ( .A0(n13712), .A1(n13746), .S(n3341), .Z(N8672) );
  CMX2X1 U24493 ( .A0(N7872), .A1(N7871), .S(n3874), .Z(n13719) );
  CMXI2X1 U24494 ( .A0(n13719), .A1(n13713), .S(n4178), .Z(n13726) );
  CMX2X1 U24495 ( .A0(n13714), .A1(n13726), .S(n3773), .Z(n13749) );
  CMXI2X1 U24496 ( .A0(n13715), .A1(n13749), .S(n3341), .Z(N8673) );
  CMX2X1 U24497 ( .A0(N7871), .A1(N7870), .S(n3875), .Z(n13722) );
  CMXI2X1 U24498 ( .A0(n13722), .A1(n13716), .S(n4178), .Z(n13729) );
  CMX2X1 U24499 ( .A0(n13717), .A1(n13729), .S(n3771), .Z(n13752) );
  CMXI2X1 U24500 ( .A0(n13718), .A1(n13752), .S(n3340), .Z(N8674) );
  CMX2X1 U24501 ( .A0(N7870), .A1(N7869), .S(n3876), .Z(n13725) );
  CMXI2X1 U24502 ( .A0(n13725), .A1(n13719), .S(n4178), .Z(n13732) );
  CMX2X1 U24503 ( .A0(n13720), .A1(n13732), .S(n3806), .Z(n13755) );
  CMXI2X1 U24504 ( .A0(n13721), .A1(n13755), .S(n3340), .Z(N8675) );
  CMX2X1 U24505 ( .A0(N7869), .A1(N7868), .S(n3877), .Z(n13728) );
  CMXI2X1 U24506 ( .A0(n13728), .A1(n13722), .S(n4178), .Z(n13745) );
  CMX2X1 U24507 ( .A0(n13723), .A1(n13745), .S(n3772), .Z(n13758) );
  CMXI2X1 U24508 ( .A0(n13724), .A1(n13758), .S(n3340), .Z(N8676) );
  CMX2X1 U24509 ( .A0(N7868), .A1(N7867), .S(n3878), .Z(n13731) );
  CMXI2X1 U24510 ( .A0(n13731), .A1(n13725), .S(n4178), .Z(n13748) );
  CMX2X1 U24511 ( .A0(n13726), .A1(n13748), .S(n3773), .Z(n13761) );
  CMXI2X1 U24512 ( .A0(n13727), .A1(n13761), .S(n3340), .Z(N8677) );
  CMX2X1 U24513 ( .A0(N7867), .A1(N7866), .S(n3879), .Z(n13744) );
  CMXI2X1 U24514 ( .A0(n13744), .A1(n13728), .S(n4178), .Z(n13751) );
  CMX2X1 U24515 ( .A0(n13729), .A1(n13751), .S(n3774), .Z(n13764) );
  CMXI2X1 U24516 ( .A0(n13730), .A1(n13764), .S(n3340), .Z(N8678) );
  CMX2X1 U24517 ( .A0(N7866), .A1(N7865), .S(n3878), .Z(n13747) );
  CMXI2X1 U24518 ( .A0(n13747), .A1(n13731), .S(n4178), .Z(n13754) );
  CMX2X1 U24519 ( .A0(n13732), .A1(n13754), .S(n3775), .Z(n13767) );
  CMXI2X1 U24520 ( .A0(n13733), .A1(n13767), .S(n3340), .Z(N8679) );
  CMX2X1 U24521 ( .A0(N8226), .A1(N8225), .S(n3879), .Z(n13807) );
  CMXI2X1 U24522 ( .A0(n13807), .A1(n13734), .S(n4178), .Z(n13873) );
  CMX2X1 U24523 ( .A0(n13735), .A1(n13873), .S(n3776), .Z(n14006) );
  CMXI2X1 U24524 ( .A0(n13736), .A1(n14006), .S(n3340), .Z(N8319) );
  CMXI2X1 U24525 ( .A0(n13738), .A1(n13737), .S(n4178), .Z(n15076) );
  CMXI2X1 U24526 ( .A0(n13743), .A1(n13742), .S(n3340), .Z(N8283) );
  CMX2X1 U24527 ( .A0(N7865), .A1(N7864), .S(n3881), .Z(n13750) );
  CMXI2X1 U24528 ( .A0(n13750), .A1(n13744), .S(n4177), .Z(n13757) );
  CMX2X1 U24529 ( .A0(n13745), .A1(n13757), .S(n3777), .Z(n13770) );
  CMX2X1 U24530 ( .A0(N7864), .A1(N7863), .S(n3862), .Z(n13753) );
  CMXI2X1 U24531 ( .A0(n13753), .A1(n13747), .S(n4177), .Z(n13760) );
  CMX2X1 U24532 ( .A0(n13748), .A1(n13760), .S(n3790), .Z(n13773) );
  CMXI2X1 U24533 ( .A0(n13749), .A1(n13773), .S(n3343), .Z(N8681) );
  CMX2X1 U24534 ( .A0(N7863), .A1(N7862), .S(n3863), .Z(n13756) );
  CMX2X1 U24535 ( .A0(n13751), .A1(n13763), .S(n3791), .Z(n13779) );
  CMXI2X1 U24536 ( .A0(n13752), .A1(n13779), .S(n3343), .Z(N8682) );
  CMX2X1 U24537 ( .A0(N7862), .A1(N7861), .S(n3864), .Z(n13759) );
  CMXI2X1 U24538 ( .A0(n13759), .A1(n13753), .S(n4177), .Z(n13766) );
  CMX2X1 U24539 ( .A0(n13754), .A1(n13766), .S(n3792), .Z(n13782) );
  CMXI2X1 U24540 ( .A0(n13755), .A1(n13782), .S(n3343), .Z(N8683) );
  CMX2X1 U24541 ( .A0(N7861), .A1(N7860), .S(n3879), .Z(n13762) );
  CMX2X1 U24542 ( .A0(n13757), .A1(n13769), .S(n3773), .Z(n13785) );
  CMXI2X1 U24543 ( .A0(n13758), .A1(n13785), .S(n3342), .Z(N8684) );
  CMX2X1 U24544 ( .A0(N7860), .A1(N7859), .S(n3880), .Z(n13765) );
  CMXI2X1 U24545 ( .A0(n13765), .A1(n13759), .S(n4177), .Z(n13772) );
  CMX2X1 U24546 ( .A0(n13760), .A1(n13772), .S(n3774), .Z(n13788) );
  CMXI2X1 U24547 ( .A0(n13761), .A1(n13788), .S(n3342), .Z(N8685) );
  CMX2X1 U24548 ( .A0(N7859), .A1(N7858), .S(n3881), .Z(n13768) );
  CMXI2X1 U24549 ( .A0(n13768), .A1(n13762), .S(n4177), .Z(n13778) );
  CMX2X1 U24550 ( .A0(n13763), .A1(n13778), .S(n3775), .Z(n13791) );
  CMXI2X1 U24551 ( .A0(n13764), .A1(n13791), .S(n3342), .Z(N8686) );
  CMX2X1 U24552 ( .A0(N7858), .A1(N7857), .S(n3862), .Z(n13771) );
  CMX2X1 U24553 ( .A0(n13766), .A1(n13781), .S(n3776), .Z(n13794) );
  CMXI2X1 U24554 ( .A0(n13767), .A1(n13794), .S(n3342), .Z(N8687) );
  CMX2X1 U24555 ( .A0(N7857), .A1(N7856), .S(n3876), .Z(n13777) );
  CMXI2X1 U24556 ( .A0(n13777), .A1(n13768), .S(n4177), .Z(n13784) );
  CMX2X1 U24557 ( .A0(n13769), .A1(n13784), .S(n3777), .Z(n13797) );
  CMXI2X1 U24558 ( .A0(n13770), .A1(n13797), .S(n3342), .Z(N8688) );
  CMX2X1 U24559 ( .A0(N7856), .A1(N7855), .S(n3880), .Z(n13780) );
  CMXI2X1 U24560 ( .A0(n13780), .A1(n13771), .S(n4177), .Z(n13787) );
  CMXI2X1 U24561 ( .A0(n13773), .A1(n13800), .S(n3342), .Z(N8689) );
  CMX2X1 U24562 ( .A0(N8225), .A1(N8224), .S(n3881), .Z(n13840) );
  CMXI2X1 U24563 ( .A0(n13840), .A1(n13774), .S(n4177), .Z(n13906) );
  CMX2X1 U24564 ( .A0(n13775), .A1(n13906), .S(n3791), .Z(n14039) );
  CMXI2X1 U24565 ( .A0(n13776), .A1(n14039), .S(n3342), .Z(N8320) );
  CMX2X1 U24566 ( .A0(N7855), .A1(N7854), .S(n3862), .Z(n13783) );
  CMXI2X1 U24567 ( .A0(n13783), .A1(n13777), .S(n4177), .Z(n13790) );
  CMX2X1 U24568 ( .A0(n13778), .A1(n13790), .S(n3776), .Z(n13803) );
  CMXI2X1 U24569 ( .A0(n13779), .A1(n13803), .S(n3342), .Z(N8690) );
  CMX2X1 U24570 ( .A0(N7854), .A1(N7853), .S(n3863), .Z(n13786) );
  CMXI2X1 U24571 ( .A0(n13786), .A1(n13780), .S(n4177), .Z(n13793) );
  CMX2X1 U24572 ( .A0(n13781), .A1(n13793), .S(n3811), .Z(n13806) );
  CMXI2X1 U24573 ( .A0(n13782), .A1(n13806), .S(n3342), .Z(N8691) );
  CMX2X1 U24574 ( .A0(N7853), .A1(N7852), .S(n3864), .Z(n13789) );
  CMXI2X1 U24575 ( .A0(n13789), .A1(n13783), .S(n4177), .Z(n13796) );
  CMX2X1 U24576 ( .A0(n13784), .A1(n13796), .S(n3808), .Z(n13812) );
  CMXI2X1 U24577 ( .A0(n13785), .A1(n13812), .S(n3342), .Z(N8692) );
  CMX2X1 U24578 ( .A0(N7852), .A1(N7851), .S(n3865), .Z(n13792) );
  CMX2X1 U24579 ( .A0(n13787), .A1(n13799), .S(n3809), .Z(n13815) );
  CMX2X1 U24580 ( .A0(N7851), .A1(N7850), .S(n3866), .Z(n13795) );
  CMXI2X1 U24581 ( .A0(n13795), .A1(n13789), .S(n4177), .Z(n13802) );
  CMX2X1 U24582 ( .A0(n13790), .A1(n13802), .S(n3810), .Z(n13818) );
  CMXI2X1 U24583 ( .A0(n13791), .A1(n13818), .S(n3342), .Z(N8694) );
  CMX2X1 U24584 ( .A0(N7850), .A1(N7849), .S(n3880), .Z(n13798) );
  CMXI2X1 U24585 ( .A0(n13798), .A1(n13792), .S(n4176), .Z(n13805) );
  CMX2X1 U24586 ( .A0(n13793), .A1(n13805), .S(n3811), .Z(n13821) );
  CMXI2X1 U24587 ( .A0(n13794), .A1(n13821), .S(n3341), .Z(N8695) );
  CMX2X1 U24588 ( .A0(N7849), .A1(N7848), .S(n3879), .Z(n13801) );
  CMXI2X1 U24589 ( .A0(n13801), .A1(n13795), .S(n4176), .Z(n13811) );
  CMX2X1 U24590 ( .A0(n13796), .A1(n13811), .S(n3812), .Z(n13824) );
  CMXI2X1 U24591 ( .A0(n13797), .A1(n13824), .S(n3341), .Z(N8696) );
  CMX2X1 U24592 ( .A0(N7848), .A1(N7847), .S(n3880), .Z(n13804) );
  CMX2X1 U24593 ( .A0(n13799), .A1(n13814), .S(n3795), .Z(n13827) );
  CMXI2X1 U24594 ( .A0(n13800), .A1(n13827), .S(n3341), .Z(N8697) );
  CMX2X1 U24595 ( .A0(N7847), .A1(N7846), .S(n3881), .Z(n13810) );
  CMXI2X1 U24596 ( .A0(n13810), .A1(n13801), .S(n4176), .Z(n13817) );
  CMX2X1 U24597 ( .A0(n13802), .A1(n13817), .S(n3792), .Z(n13830) );
  CMXI2X1 U24598 ( .A0(n13803), .A1(n13830), .S(n3344), .Z(N8698) );
  CMX2X1 U24599 ( .A0(N7846), .A1(N7845), .S(n3865), .Z(n13813) );
  CMXI2X1 U24600 ( .A0(n13813), .A1(n13804), .S(n4176), .Z(n13820) );
  CMX2X1 U24601 ( .A0(n13805), .A1(n13820), .S(n3793), .Z(n13833) );
  CMXI2X1 U24602 ( .A0(n13806), .A1(n13833), .S(n3344), .Z(N8699) );
  CMX2X1 U24603 ( .A0(N8224), .A1(N8223), .S(n3875), .Z(n13872) );
  CMXI2X1 U24604 ( .A0(n13872), .A1(n13807), .S(n4176), .Z(n13939) );
  CMX2X1 U24605 ( .A0(n13808), .A1(n13939), .S(n3794), .Z(n14072) );
  CMXI2X1 U24606 ( .A0(n13809), .A1(n14072), .S(n3344), .Z(N8321) );
  CMX2X1 U24607 ( .A0(N7845), .A1(N7844), .S(n3876), .Z(n13816) );
  CMXI2X1 U24608 ( .A0(n13816), .A1(n13810), .S(n4176), .Z(n13823) );
  CMX2X1 U24609 ( .A0(n13811), .A1(n13823), .S(n3795), .Z(n13836) );
  CMXI2X1 U24610 ( .A0(n13812), .A1(n13836), .S(n3344), .Z(N8700) );
  CMX2X1 U24611 ( .A0(N7844), .A1(N7843), .S(n3877), .Z(n13819) );
  CMXI2X1 U24612 ( .A0(n13819), .A1(n13813), .S(n4176), .Z(n13826) );
  CMX2X1 U24613 ( .A0(n13814), .A1(n13826), .S(n3796), .Z(n13839) );
  CMXI2X1 U24614 ( .A0(n13815), .A1(n13839), .S(n3344), .Z(N8701) );
  CMX2X1 U24615 ( .A0(N7843), .A1(N7842), .S(n3878), .Z(n13822) );
  CMXI2X1 U24616 ( .A0(n13822), .A1(n13816), .S(n4176), .Z(n13829) );
  CMX2X1 U24617 ( .A0(n13817), .A1(n13829), .S(n3797), .Z(n13845) );
  CMXI2X1 U24618 ( .A0(n13818), .A1(n13845), .S(n3344), .Z(N8702) );
  CMX2X1 U24619 ( .A0(N7842), .A1(N7841), .S(n3879), .Z(n13825) );
  CMX2X1 U24620 ( .A0(n13820), .A1(n13832), .S(n3805), .Z(n13848) );
  CMXI2X1 U24621 ( .A0(n13821), .A1(n13848), .S(n3344), .Z(N8703) );
  CMX2X1 U24622 ( .A0(N7841), .A1(N7840), .S(n3880), .Z(n13828) );
  CMXI2X1 U24623 ( .A0(n13828), .A1(n13822), .S(n4176), .Z(n13835) );
  CMX2X1 U24624 ( .A0(n13823), .A1(n13835), .S(n3806), .Z(n13851) );
  CMXI2X1 U24625 ( .A0(n13824), .A1(n13851), .S(n3344), .Z(N8704) );
  CMX2X1 U24626 ( .A0(N7840), .A1(N7839), .S(n3881), .Z(n13831) );
  CMXI2X1 U24627 ( .A0(n13831), .A1(n13825), .S(n4176), .Z(n13838) );
  CMX2X1 U24628 ( .A0(n13826), .A1(n13838), .S(n3807), .Z(n13854) );
  CMXI2X1 U24629 ( .A0(n13827), .A1(n13854), .S(n3344), .Z(N8705) );
  CMX2X1 U24630 ( .A0(N7839), .A1(N7838), .S(n3869), .Z(n13834) );
  CMXI2X1 U24631 ( .A0(n13834), .A1(n13828), .S(n4176), .Z(n13844) );
  CMX2X1 U24632 ( .A0(n13829), .A1(n13844), .S(n3808), .Z(n13857) );
  CMXI2X1 U24633 ( .A0(n13830), .A1(n13857), .S(n3343), .Z(N8706) );
  CMX2X1 U24634 ( .A0(N7838), .A1(N7837), .S(n3870), .Z(n13837) );
  CMX2X1 U24635 ( .A0(n13832), .A1(n13847), .S(n3809), .Z(n13859) );
  CMXI2X1 U24636 ( .A0(n13833), .A1(n13859), .S(n3343), .Z(N8707) );
  CMX2X1 U24637 ( .A0(N7837), .A1(N7836), .S(n3862), .Z(n13843) );
  CMXI2X1 U24638 ( .A0(n13843), .A1(n13834), .S(n4176), .Z(n13850) );
  CMX2X1 U24639 ( .A0(n13835), .A1(n13850), .S(n3810), .Z(n13862) );
  CMXI2X1 U24640 ( .A0(n13836), .A1(n13862), .S(n3343), .Z(N8708) );
  CMX2X1 U24641 ( .A0(N7836), .A1(N7835), .S(n3863), .Z(n13846) );
  CMXI2X1 U24642 ( .A0(n13846), .A1(n13837), .S(n4176), .Z(n13853) );
  CMX2X1 U24643 ( .A0(n13838), .A1(n13853), .S(n3811), .Z(n13865) );
  CMXI2X1 U24644 ( .A0(n13839), .A1(n13865), .S(n3343), .Z(N8709) );
  CMX2X1 U24645 ( .A0(N8223), .A1(N8222), .S(n3869), .Z(n13905) );
  CMXI2X1 U24646 ( .A0(n13905), .A1(n13840), .S(n4175), .Z(n13972) );
  CMX2X1 U24647 ( .A0(n13841), .A1(n13972), .S(n3812), .Z(n14109) );
  CMXI2X1 U24648 ( .A0(n13842), .A1(n14109), .S(n3343), .Z(N8322) );
  CMX2X1 U24649 ( .A0(N7835), .A1(N7834), .S(n3870), .Z(n13849) );
  CMX2X1 U24650 ( .A0(n13844), .A1(n13856), .S(n4365), .Z(n13868) );
  CMX2X1 U24651 ( .A0(N7834), .A1(N7833), .S(n3871), .Z(n13852) );
  CMX2X1 U24652 ( .A0(n13847), .A1(n13858), .S(n3771), .Z(n13871) );
  CMX2X1 U24653 ( .A0(N7833), .A1(N7832), .S(n3872), .Z(n13855) );
  CMXI2X1 U24654 ( .A0(n13855), .A1(n13849), .S(n4175), .Z(n13861) );
  CMX2X1 U24655 ( .A0(n13850), .A1(n13861), .S(n3777), .Z(n13877) );
  CMXI2X1 U24656 ( .A0(n13851), .A1(n13877), .S(n3343), .Z(N8712) );
  CMX2X1 U24657 ( .A0(n13853), .A1(n13864), .S(n3812), .Z(n13880) );
  CMX2X1 U24658 ( .A0(N7831), .A1(N7830), .S(n3863), .Z(n13860) );
  CMXI2X1 U24659 ( .A0(n13860), .A1(n13855), .S(n4175), .Z(n13867) );
  CMX2X1 U24660 ( .A0(n13856), .A1(n13867), .S(n4368), .Z(n13883) );
  CMXI2X1 U24661 ( .A0(n13857), .A1(n13883), .S(n3346), .Z(N8714) );
  CMX2X1 U24662 ( .A0(N7830), .A1(N7829), .S(n3864), .Z(n13863) );
  CMXI2X1 U24663 ( .A0(n13863), .A1(n3707), .S(n4175), .Z(n13870) );
  CMX2X1 U24664 ( .A0(n3704), .A1(n13870), .S(n3771), .Z(n13886) );
  CMXI2X1 U24665 ( .A0(n13859), .A1(n13886), .S(n3345), .Z(N8715) );
  CMX2X1 U24666 ( .A0(N7829), .A1(N7828), .S(n3881), .Z(n13866) );
  CMXI2X1 U24667 ( .A0(n13866), .A1(n13860), .S(n4175), .Z(n13876) );
  CMX2X1 U24668 ( .A0(n13861), .A1(n13876), .S(n3772), .Z(n13889) );
  CMXI2X1 U24669 ( .A0(n13862), .A1(n13889), .S(n3345), .Z(N8716) );
  CMX2X1 U24670 ( .A0(N7828), .A1(N7827), .S(n3867), .Z(n13869) );
  CMXI2X1 U24671 ( .A0(n13869), .A1(n13863), .S(n4175), .Z(n13879) );
  CMX2X1 U24672 ( .A0(n13864), .A1(n13879), .S(n3773), .Z(n13892) );
  CMXI2X1 U24673 ( .A0(n13865), .A1(n13892), .S(n3345), .Z(N8717) );
  CMX2X1 U24674 ( .A0(N7827), .A1(N7826), .S(n3868), .Z(n13875) );
  CMXI2X1 U24675 ( .A0(n13875), .A1(n13866), .S(n4175), .Z(n13882) );
  CMX2X1 U24676 ( .A0(n13867), .A1(n13882), .S(n3774), .Z(n13895) );
  CMXI2X1 U24677 ( .A0(n13868), .A1(n13895), .S(n3345), .Z(N8718) );
  CMX2X1 U24678 ( .A0(N7826), .A1(N7825), .S(n3865), .Z(n13878) );
  CMXI2X1 U24679 ( .A0(n13878), .A1(n13869), .S(n4175), .Z(n13885) );
  CMX2X1 U24680 ( .A0(n13870), .A1(n13885), .S(n3796), .Z(n13898) );
  CMXI2X1 U24681 ( .A0(n13871), .A1(n13898), .S(n3345), .Z(N8719) );
  CMX2X1 U24682 ( .A0(N8222), .A1(N8221), .S(n3866), .Z(n13938) );
  CMXI2X1 U24683 ( .A0(n13938), .A1(n13872), .S(n4175), .Z(n14005) );
  CMX2X1 U24684 ( .A0(n13873), .A1(n14005), .S(n3772), .Z(n14142) );
  CMXI2X1 U24685 ( .A0(n13874), .A1(n14142), .S(n3345), .Z(N8323) );
  CMX2X1 U24686 ( .A0(N7825), .A1(N7824), .S(n3867), .Z(n13881) );
  CMXI2X1 U24687 ( .A0(n13881), .A1(n13875), .S(n4175), .Z(n13888) );
  CMX2X1 U24688 ( .A0(n13876), .A1(n13888), .S(n3773), .Z(n13901) );
  CMX2X1 U24689 ( .A0(N7824), .A1(N7823), .S(n3868), .Z(n13884) );
  CMXI2X1 U24690 ( .A0(n13884), .A1(n13878), .S(n4175), .Z(n13891) );
  CMX2X1 U24691 ( .A0(n13879), .A1(n13891), .S(n3774), .Z(n13904) );
  CMXI2X1 U24692 ( .A0(n13880), .A1(n13904), .S(n3345), .Z(N8721) );
  CMX2X1 U24693 ( .A0(N7823), .A1(N7822), .S(n3863), .Z(n13887) );
  CMXI2X1 U24694 ( .A0(n13887), .A1(n13881), .S(n4175), .Z(n13894) );
  CMX2X1 U24695 ( .A0(n13882), .A1(n13894), .S(n3775), .Z(n13910) );
  CMX2X1 U24696 ( .A0(N7822), .A1(N7821), .S(n3864), .Z(n13890) );
  CMXI2X1 U24697 ( .A0(n13890), .A1(n13884), .S(n4175), .Z(n13897) );
  CMX2X1 U24698 ( .A0(n13885), .A1(n13897), .S(n3776), .Z(n13913) );
  CMXI2X1 U24699 ( .A0(n13886), .A1(n13913), .S(n3345), .Z(N8723) );
  CMX2X1 U24700 ( .A0(N7821), .A1(N7820), .S(n3865), .Z(n13893) );
  CMXI2X1 U24701 ( .A0(n13893), .A1(n13887), .S(n4174), .Z(n13900) );
  CMX2X1 U24702 ( .A0(n13888), .A1(n13900), .S(n3777), .Z(n13916) );
  CMX2X1 U24703 ( .A0(N7820), .A1(N7819), .S(n3866), .Z(n13896) );
  CMX2X1 U24704 ( .A0(n13891), .A1(n13903), .S(n3790), .Z(n13919) );
  CMXI2X1 U24705 ( .A0(n13892), .A1(n13919), .S(n3345), .Z(N8725) );
  CMX2X1 U24706 ( .A0(N7819), .A1(N7818), .S(n3877), .Z(n13899) );
  CMXI2X1 U24707 ( .A0(n13899), .A1(n13893), .S(n4174), .Z(n13909) );
  CMX2X1 U24708 ( .A0(n13894), .A1(n13909), .S(n3791), .Z(n13922) );
  CMXI2X1 U24709 ( .A0(n13895), .A1(n13922), .S(n3345), .Z(N8726) );
  CMX2X1 U24710 ( .A0(N7818), .A1(N7817), .S(n3869), .Z(n13902) );
  CMXI2X1 U24711 ( .A0(n13902), .A1(n13896), .S(n4174), .Z(n13912) );
  CMX2X1 U24712 ( .A0(n13897), .A1(n13912), .S(n3792), .Z(n13925) );
  CMXI2X1 U24713 ( .A0(n13898), .A1(n13925), .S(n3345), .Z(N8727) );
  CMX2X1 U24714 ( .A0(N7817), .A1(N7816), .S(n3870), .Z(n13908) );
  CMXI2X1 U24715 ( .A0(n13908), .A1(n13899), .S(n4174), .Z(n13915) );
  CMX2X1 U24716 ( .A0(n13900), .A1(n13915), .S(n3793), .Z(n13928) );
  CMXI2X1 U24717 ( .A0(n13901), .A1(n13928), .S(n3344), .Z(N8728) );
  CMX2X1 U24718 ( .A0(N7816), .A1(N7815), .S(n3871), .Z(n13911) );
  CMXI2X1 U24719 ( .A0(n13911), .A1(n13902), .S(n4174), .Z(n13918) );
  CMX2X1 U24720 ( .A0(n13903), .A1(n13918), .S(n3794), .Z(n13931) );
  CMXI2X1 U24721 ( .A0(n13904), .A1(n13931), .S(n3344), .Z(N8729) );
  CMX2X1 U24722 ( .A0(N8221), .A1(N8220), .S(n3872), .Z(n13971) );
  CMXI2X1 U24723 ( .A0(n13971), .A1(n13905), .S(n4174), .Z(n14038) );
  CMX2X1 U24724 ( .A0(n13906), .A1(n14038), .S(n3795), .Z(n14175) );
  CMX2X1 U24725 ( .A0(N7815), .A1(N7814), .S(n3873), .Z(n13914) );
  CMXI2X1 U24726 ( .A0(n13914), .A1(n13908), .S(n4174), .Z(n13921) );
  CMX2X1 U24727 ( .A0(n13909), .A1(n13921), .S(n3796), .Z(n13934) );
  CMXI2X1 U24728 ( .A0(n13910), .A1(n13934), .S(n3347), .Z(N8730) );
  CMX2X1 U24729 ( .A0(N7814), .A1(N7813), .S(n3874), .Z(n13917) );
  CMXI2X1 U24730 ( .A0(n13917), .A1(n13911), .S(n4174), .Z(n13924) );
  CMX2X1 U24731 ( .A0(n13912), .A1(n13924), .S(n3797), .Z(n13937) );
  CMXI2X1 U24732 ( .A0(n13913), .A1(n13937), .S(n3347), .Z(N8731) );
  CMX2X1 U24733 ( .A0(N7813), .A1(N7812), .S(n3875), .Z(n13920) );
  CMX2X1 U24734 ( .A0(n13915), .A1(n13927), .S(n3805), .Z(n13943) );
  CMXI2X1 U24735 ( .A0(n13916), .A1(n13943), .S(n3347), .Z(N8732) );
  CMX2X1 U24736 ( .A0(N7812), .A1(N7811), .S(n3862), .Z(n13923) );
  CMX2X1 U24737 ( .A0(n13918), .A1(n13930), .S(n3806), .Z(n13946) );
  CMXI2X1 U24738 ( .A0(n13919), .A1(n13946), .S(n3347), .Z(N8733) );
  CMX2X1 U24739 ( .A0(N7811), .A1(N7810), .S(n3871), .Z(n13926) );
  CMXI2X1 U24740 ( .A0(n13926), .A1(n13920), .S(n4174), .Z(n13933) );
  CMX2X1 U24741 ( .A0(n13921), .A1(n13933), .S(n3790), .Z(n13949) );
  CMXI2X1 U24742 ( .A0(n13922), .A1(n13949), .S(n3347), .Z(N8734) );
  CMX2X1 U24743 ( .A0(N7810), .A1(N7809), .S(n3868), .Z(n13929) );
  CMXI2X1 U24744 ( .A0(n13929), .A1(n13923), .S(n4174), .Z(n13936) );
  CMX2X1 U24745 ( .A0(n13924), .A1(n13936), .S(n4306), .Z(n13952) );
  CMXI2X1 U24746 ( .A0(n13925), .A1(n13952), .S(n3347), .Z(N8735) );
  CMX2X1 U24747 ( .A0(N7809), .A1(N7808), .S(n3863), .Z(n13932) );
  CMXI2X1 U24748 ( .A0(n13932), .A1(n13926), .S(n4174), .Z(n13942) );
  CMX2X1 U24749 ( .A0(n13927), .A1(n13942), .S(n3775), .Z(n13955) );
  CMXI2X1 U24750 ( .A0(n13928), .A1(n13955), .S(n3347), .Z(N8736) );
  CMX2X1 U24751 ( .A0(N7808), .A1(N7807), .S(n3864), .Z(n13935) );
  CMXI2X1 U24752 ( .A0(n13935), .A1(n13929), .S(n4174), .Z(n13945) );
  CMX2X1 U24753 ( .A0(n13930), .A1(n13945), .S(n3776), .Z(n13958) );
  CMXI2X1 U24754 ( .A0(n13931), .A1(n13958), .S(n3347), .Z(N8737) );
  CMX2X1 U24755 ( .A0(N7807), .A1(N7806), .S(n3865), .Z(n13941) );
  CMXI2X1 U24756 ( .A0(n13941), .A1(n13932), .S(n4174), .Z(n13948) );
  CMX2X1 U24757 ( .A0(n13933), .A1(n13948), .S(n3777), .Z(n13961) );
  CMXI2X1 U24758 ( .A0(n13934), .A1(n13961), .S(n3346), .Z(N8738) );
  CMX2X1 U24759 ( .A0(N7806), .A1(N7805), .S(n3866), .Z(n13944) );
  CMXI2X1 U24760 ( .A0(n13944), .A1(n13935), .S(n4173), .Z(n13951) );
  CMX2X1 U24761 ( .A0(n13936), .A1(n13951), .S(n3790), .Z(n13964) );
  CMXI2X1 U24762 ( .A0(n13937), .A1(n13964), .S(n3346), .Z(N8739) );
  CMX2X1 U24763 ( .A0(N8220), .A1(N8219), .S(n3862), .Z(n14004) );
  CMXI2X1 U24764 ( .A0(n14004), .A1(n13938), .S(n4173), .Z(n14071) );
  CMX2X1 U24765 ( .A0(n13939), .A1(n14071), .S(n3791), .Z(n14208) );
  CMXI2X1 U24766 ( .A0(n13940), .A1(n14208), .S(n3346), .Z(N8325) );
  CMX2X1 U24767 ( .A0(N7805), .A1(N7804), .S(n3874), .Z(n13947) );
  CMXI2X1 U24768 ( .A0(n13947), .A1(n13941), .S(n4173), .Z(n13954) );
  CMX2X1 U24769 ( .A0(n13942), .A1(n13954), .S(n3797), .Z(n13967) );
  CMXI2X1 U24770 ( .A0(n13943), .A1(n13967), .S(n3346), .Z(N8740) );
  CMX2X1 U24771 ( .A0(N7804), .A1(N7803), .S(n3875), .Z(n13950) );
  CMXI2X1 U24772 ( .A0(n13950), .A1(n13944), .S(n4173), .Z(n13957) );
  CMX2X1 U24773 ( .A0(n13945), .A1(n13957), .S(n3807), .Z(n13970) );
  CMXI2X1 U24774 ( .A0(n13946), .A1(n13970), .S(n3346), .Z(N8741) );
  CMX2X1 U24775 ( .A0(N7803), .A1(N7802), .S(n3876), .Z(n13953) );
  CMXI2X1 U24776 ( .A0(n13953), .A1(n13947), .S(n4173), .Z(n13960) );
  CMX2X1 U24777 ( .A0(n13948), .A1(n13960), .S(n3808), .Z(n13976) );
  CMXI2X1 U24778 ( .A0(n13949), .A1(n13976), .S(n3346), .Z(N8742) );
  CMX2X1 U24779 ( .A0(N7802), .A1(N7801), .S(n3877), .Z(n13956) );
  CMX2X1 U24780 ( .A0(n13951), .A1(n13963), .S(n3809), .Z(n13979) );
  CMXI2X1 U24781 ( .A0(n13952), .A1(n13979), .S(n3346), .Z(N8743) );
  CMX2X1 U24782 ( .A0(N7801), .A1(N7800), .S(n3878), .Z(n13959) );
  CMXI2X1 U24783 ( .A0(n13959), .A1(n13953), .S(n4173), .Z(n13966) );
  CMX2X1 U24784 ( .A0(n13954), .A1(n13966), .S(n3810), .Z(n13982) );
  CMXI2X1 U24785 ( .A0(n13955), .A1(n13982), .S(n3346), .Z(N8744) );
  CMX2X1 U24786 ( .A0(N7800), .A1(N7799), .S(n3879), .Z(n13962) );
  CMXI2X1 U24787 ( .A0(n13962), .A1(n13956), .S(n4173), .Z(n13969) );
  CMX2X1 U24788 ( .A0(n13957), .A1(n13969), .S(n3811), .Z(n13985) );
  CMXI2X1 U24789 ( .A0(n13958), .A1(n13985), .S(n3346), .Z(N8745) );
  CMX2X1 U24790 ( .A0(N7799), .A1(N7798), .S(n3880), .Z(n13965) );
  CMXI2X1 U24791 ( .A0(n13965), .A1(n13959), .S(n4173), .Z(n13975) );
  CMX2X1 U24792 ( .A0(n13960), .A1(n13975), .S(n3812), .Z(n13988) );
  CMXI2X1 U24793 ( .A0(n13961), .A1(n13988), .S(n3346), .Z(N8746) );
  CMX2X1 U24794 ( .A0(N7798), .A1(N7797), .S(n3872), .Z(n13968) );
  CMXI2X1 U24795 ( .A0(n13968), .A1(n13962), .S(n4173), .Z(n13978) );
  CMX2X1 U24796 ( .A0(n13963), .A1(n13978), .S(n4305), .Z(n13991) );
  CMXI2X1 U24797 ( .A0(n13964), .A1(n13991), .S(n3496), .Z(N8747) );
  CMX2X1 U24798 ( .A0(N7797), .A1(N7796), .S(n3873), .Z(n13974) );
  CMXI2X1 U24799 ( .A0(n13974), .A1(n13965), .S(n4173), .Z(n13981) );
  CMX2X1 U24800 ( .A0(n13966), .A1(n13981), .S(n3811), .Z(n13994) );
  CMXI2X1 U24801 ( .A0(n13967), .A1(n13994), .S(n3495), .Z(N8748) );
  CMX2X1 U24802 ( .A0(N7796), .A1(N7795), .S(n3881), .Z(n13977) );
  CMXI2X1 U24803 ( .A0(n13977), .A1(n13968), .S(n4173), .Z(n13984) );
  CMX2X1 U24804 ( .A0(n13969), .A1(n13984), .S(n4322), .Z(n13997) );
  CMXI2X1 U24805 ( .A0(n13970), .A1(n13997), .S(n3494), .Z(N8749) );
  CMX2X1 U24806 ( .A0(N8219), .A1(N8218), .S(n3862), .Z(n14037) );
  CMX2X1 U24807 ( .A0(n13972), .A1(n14108), .S(n4321), .Z(n14241) );
  CMXI2X1 U24808 ( .A0(n13973), .A1(n14241), .S(n3386), .Z(N8326) );
  CMX2X1 U24809 ( .A0(N7795), .A1(N7794), .S(n3869), .Z(n13980) );
  CMXI2X1 U24810 ( .A0(n13980), .A1(n13974), .S(n4173), .Z(n13987) );
  CMX2X1 U24811 ( .A0(n13975), .A1(n13987), .S(n4321), .Z(n14000) );
  CMXI2X1 U24812 ( .A0(n13976), .A1(n14000), .S(n3348), .Z(N8750) );
  CMX2X1 U24813 ( .A0(N7794), .A1(N7793), .S(n3870), .Z(n13983) );
  CMX2X1 U24814 ( .A0(n13978), .A1(n13990), .S(n4321), .Z(n14003) );
  CMXI2X1 U24815 ( .A0(n13979), .A1(n14003), .S(n3348), .Z(N8751) );
  CMX2X1 U24816 ( .A0(N7793), .A1(N7792), .S(n3871), .Z(n13986) );
  CMXI2X1 U24817 ( .A0(n13986), .A1(n13980), .S(n4173), .Z(n13993) );
  CMX2X1 U24818 ( .A0(n13981), .A1(n13993), .S(n4321), .Z(n14009) );
  CMXI2X1 U24819 ( .A0(n13982), .A1(n14009), .S(n3348), .Z(N8752) );
  CMX2X1 U24820 ( .A0(N7792), .A1(N7791), .S(n3872), .Z(n13989) );
  CMXI2X1 U24821 ( .A0(n13989), .A1(n13983), .S(n4172), .Z(n13996) );
  CMX2X1 U24822 ( .A0(n13984), .A1(n13996), .S(n4321), .Z(n14012) );
  CMXI2X1 U24823 ( .A0(n13985), .A1(n14012), .S(n3348), .Z(N8753) );
  CMX2X1 U24824 ( .A0(N7791), .A1(N7790), .S(n3867), .Z(n13992) );
  CMXI2X1 U24825 ( .A0(n13992), .A1(n13986), .S(n4172), .Z(n13999) );
  CMX2X1 U24826 ( .A0(n13987), .A1(n13999), .S(n4321), .Z(n14015) );
  CMXI2X1 U24827 ( .A0(n13988), .A1(n14015), .S(n3348), .Z(N8754) );
  CMX2X1 U24828 ( .A0(N7790), .A1(N7789), .S(n3868), .Z(n13995) );
  CMXI2X1 U24829 ( .A0(n13995), .A1(n13989), .S(n4172), .Z(n14002) );
  CMX2X1 U24830 ( .A0(n13990), .A1(n14002), .S(n4321), .Z(n14018) );
  CMXI2X1 U24831 ( .A0(n13991), .A1(n14018), .S(n3348), .Z(N8755) );
  CMXI2X1 U24832 ( .A0(n13998), .A1(n13992), .S(n4172), .Z(n14008) );
  CMX2X1 U24833 ( .A0(n13993), .A1(n14008), .S(n4321), .Z(n14021) );
  CMXI2X1 U24834 ( .A0(n13994), .A1(n14021), .S(n3348), .Z(N8756) );
  CMX2X1 U24835 ( .A0(N7788), .A1(N7787), .S(n3870), .Z(n14001) );
  CMX2X1 U24836 ( .A0(n13996), .A1(n14011), .S(n4321), .Z(n14024) );
  CMXI2X1 U24837 ( .A0(n13997), .A1(n14024), .S(n3348), .Z(N8757) );
  CMX2X1 U24838 ( .A0(N7787), .A1(N7786), .S(n3863), .Z(n14007) );
  CMX2X1 U24839 ( .A0(n13999), .A1(n14014), .S(n4321), .Z(n14027) );
  CMXI2X1 U24840 ( .A0(n14000), .A1(n14027), .S(n3348), .Z(N8758) );
  CMX2X1 U24841 ( .A0(N7786), .A1(N7785), .S(n3863), .Z(n14010) );
  CMX2X1 U24842 ( .A0(n14002), .A1(n14017), .S(n4321), .Z(n14030) );
  CMXI2X1 U24843 ( .A0(n14003), .A1(n14030), .S(n3348), .Z(N8759) );
  CMX2X1 U24844 ( .A0(N8218), .A1(N8217), .S(n3864), .Z(n14070) );
  CMXI2X1 U24845 ( .A0(n14070), .A1(n14004), .S(n4172), .Z(n14141) );
  CMX2X1 U24846 ( .A0(n14005), .A1(n14141), .S(n4320), .Z(n14274) );
  CMXI2X1 U24847 ( .A0(n14006), .A1(n14274), .S(n3348), .Z(N8327) );
  CMX2X1 U24848 ( .A0(N7785), .A1(N7784), .S(n3865), .Z(n14013) );
  CMX2X1 U24849 ( .A0(n14008), .A1(n14020), .S(n4320), .Z(n14033) );
  CMXI2X1 U24850 ( .A0(n14009), .A1(n14033), .S(n3347), .Z(N8760) );
  CMX2X1 U24851 ( .A0(N7784), .A1(N7783), .S(n3866), .Z(n14016) );
  CMXI2X1 U24852 ( .A0(n14016), .A1(n14010), .S(n4172), .Z(n14023) );
  CMX2X1 U24853 ( .A0(n14011), .A1(n14023), .S(n4320), .Z(n14036) );
  CMXI2X1 U24854 ( .A0(n14012), .A1(n14036), .S(n3347), .Z(N8761) );
  CMX2X1 U24855 ( .A0(N7783), .A1(N7782), .S(n3867), .Z(n14019) );
  CMXI2X1 U24856 ( .A0(n14019), .A1(n14013), .S(n4172), .Z(n14026) );
  CMX2X1 U24857 ( .A0(n14014), .A1(n14026), .S(n4320), .Z(n14042) );
  CMXI2X1 U24858 ( .A0(n14015), .A1(n14042), .S(n3356), .Z(N8762) );
  CMX2X1 U24859 ( .A0(N7782), .A1(N7781), .S(n3868), .Z(n14022) );
  CMXI2X1 U24860 ( .A0(n14022), .A1(n14016), .S(n4172), .Z(n14029) );
  CMX2X1 U24861 ( .A0(n14017), .A1(n14029), .S(n4320), .Z(n14045) );
  CMXI2X1 U24862 ( .A0(n14018), .A1(n14045), .S(n3349), .Z(N8763) );
  CMX2X1 U24863 ( .A0(N7781), .A1(N7780), .S(n3869), .Z(n14025) );
  CMXI2X1 U24864 ( .A0(n14025), .A1(n14019), .S(n4172), .Z(n14032) );
  CMX2X1 U24865 ( .A0(n14020), .A1(n14032), .S(n4320), .Z(n14048) );
  CMXI2X1 U24866 ( .A0(n14021), .A1(n14048), .S(n3349), .Z(N8764) );
  CMX2X1 U24867 ( .A0(N7780), .A1(N7779), .S(n3874), .Z(n14028) );
  CMXI2X1 U24868 ( .A0(n14028), .A1(n14022), .S(n4172), .Z(n14035) );
  CMX2X1 U24869 ( .A0(n14023), .A1(n14035), .S(n4320), .Z(n14051) );
  CMXI2X1 U24870 ( .A0(n14024), .A1(n14051), .S(n3349), .Z(N8765) );
  CMX2X1 U24871 ( .A0(N7779), .A1(N7778), .S(n3875), .Z(n14031) );
  CMXI2X1 U24872 ( .A0(n14031), .A1(n14025), .S(n4172), .Z(n14041) );
  CMX2X1 U24873 ( .A0(n14026), .A1(n14041), .S(n4320), .Z(n14054) );
  CMXI2X1 U24874 ( .A0(n14027), .A1(n14054), .S(n3357), .Z(N8766) );
  CMX2X1 U24875 ( .A0(N7778), .A1(N7777), .S(n3870), .Z(n14034) );
  CMXI2X1 U24876 ( .A0(n14034), .A1(n14028), .S(n4172), .Z(n14044) );
  CMX2X1 U24877 ( .A0(n14029), .A1(n14044), .S(n4320), .Z(n14057) );
  CMX2X1 U24878 ( .A0(N7777), .A1(N7776), .S(n3871), .Z(n14040) );
  CMXI2X1 U24879 ( .A0(n14040), .A1(n14031), .S(n4171), .Z(n14047) );
  CMX2X1 U24880 ( .A0(n14032), .A1(n14047), .S(n4320), .Z(n14060) );
  CMXI2X1 U24881 ( .A0(n14033), .A1(n14060), .S(n3357), .Z(N8768) );
  CMX2X1 U24882 ( .A0(N7776), .A1(N7775), .S(n3873), .Z(n14043) );
  CMXI2X1 U24883 ( .A0(n14043), .A1(n14034), .S(n4171), .Z(n14050) );
  CMX2X1 U24884 ( .A0(n14035), .A1(n14050), .S(n4320), .Z(n14063) );
  CMXI2X1 U24885 ( .A0(n14036), .A1(n14063), .S(n3351), .Z(N8769) );
  CMX2X1 U24886 ( .A0(N8217), .A1(N8216), .S(n3874), .Z(n14107) );
  CMXI2X1 U24887 ( .A0(n14107), .A1(n14037), .S(n4171), .Z(n14174) );
  CMX2X1 U24888 ( .A0(n14038), .A1(n14174), .S(n4319), .Z(n14307) );
  CMXI2X1 U24889 ( .A0(n14039), .A1(n14307), .S(n3351), .Z(N8328) );
  CMX2X1 U24890 ( .A0(N7775), .A1(N7774), .S(n3875), .Z(n14046) );
  CMXI2X1 U24891 ( .A0(n14046), .A1(n14040), .S(n4171), .Z(n14053) );
  CMX2X1 U24892 ( .A0(n14041), .A1(n14053), .S(n4319), .Z(n14066) );
  CMXI2X1 U24893 ( .A0(n14042), .A1(n14066), .S(n3351), .Z(N8770) );
  CMX2X1 U24894 ( .A0(N7774), .A1(N7773), .S(n3876), .Z(n14049) );
  CMXI2X1 U24895 ( .A0(n14049), .A1(n14043), .S(n4171), .Z(n14056) );
  CMX2X1 U24896 ( .A0(n14044), .A1(n14056), .S(n4319), .Z(n14069) );
  CMXI2X1 U24897 ( .A0(n14045), .A1(n14069), .S(n3351), .Z(N8771) );
  CMX2X1 U24898 ( .A0(N7773), .A1(N7772), .S(n3871), .Z(n14052) );
  CMXI2X1 U24899 ( .A0(n14052), .A1(n14046), .S(n4171), .Z(n14059) );
  CMX2X1 U24900 ( .A0(n14047), .A1(n14059), .S(n4319), .Z(n14079) );
  CMXI2X1 U24901 ( .A0(n14048), .A1(n14079), .S(n3351), .Z(N8772) );
  CMX2X1 U24902 ( .A0(N7772), .A1(N7771), .S(n3872), .Z(n14055) );
  CMXI2X1 U24903 ( .A0(n14055), .A1(n14049), .S(n4171), .Z(n14062) );
  CMX2X1 U24904 ( .A0(n14050), .A1(n14062), .S(n4319), .Z(n14082) );
  CMXI2X1 U24905 ( .A0(n14051), .A1(n14082), .S(n3351), .Z(N8773) );
  CMX2X1 U24906 ( .A0(N7771), .A1(N7770), .S(n3873), .Z(n14058) );
  CMXI2X1 U24907 ( .A0(n14058), .A1(n14052), .S(n4171), .Z(n14065) );
  CMX2X1 U24908 ( .A0(n14053), .A1(n14065), .S(n4319), .Z(n14085) );
  CMXI2X1 U24909 ( .A0(n14054), .A1(n14085), .S(n3351), .Z(N8774) );
  CMX2X1 U24910 ( .A0(N7770), .A1(N7769), .S(n3874), .Z(n14061) );
  CMXI2X1 U24911 ( .A0(n14061), .A1(n14055), .S(n4171), .Z(n14068) );
  CMX2X1 U24912 ( .A0(n14056), .A1(n14068), .S(n4319), .Z(n14088) );
  CMXI2X1 U24913 ( .A0(n14057), .A1(n14088), .S(n3351), .Z(N8775) );
  CMX2X1 U24914 ( .A0(N7769), .A1(N7768), .S(n3864), .Z(n14064) );
  CMXI2X1 U24915 ( .A0(n14064), .A1(n14058), .S(n4171), .Z(n14078) );
  CMX2X1 U24916 ( .A0(n14059), .A1(n14078), .S(n4319), .Z(n14091) );
  CMXI2X1 U24917 ( .A0(n14060), .A1(n14091), .S(n3351), .Z(N8776) );
  CMX2X1 U24918 ( .A0(N7768), .A1(N7767), .S(n3872), .Z(n14067) );
  CMXI2X1 U24919 ( .A0(n14067), .A1(n14061), .S(n4171), .Z(n14081) );
  CMX2X1 U24920 ( .A0(n14062), .A1(n14081), .S(n4319), .Z(n14094) );
  CMXI2X1 U24921 ( .A0(n14063), .A1(n14094), .S(n3351), .Z(N8777) );
  CMX2X1 U24922 ( .A0(N7767), .A1(N7766), .S(n3873), .Z(n14077) );
  CMXI2X1 U24923 ( .A0(n14077), .A1(n14064), .S(n4171), .Z(n14084) );
  CMX2X1 U24924 ( .A0(n14065), .A1(n14084), .S(n4319), .Z(n14097) );
  CMXI2X1 U24925 ( .A0(n14066), .A1(n14097), .S(n3351), .Z(N8778) );
  CMX2X1 U24926 ( .A0(N7766), .A1(N7765), .S(n3874), .Z(n14080) );
  CMXI2X1 U24927 ( .A0(n14080), .A1(n14067), .S(n4171), .Z(n14087) );
  CMX2X1 U24928 ( .A0(n14068), .A1(n14087), .S(n4319), .Z(n14100) );
  CMXI2X1 U24929 ( .A0(n14069), .A1(n14100), .S(n3350), .Z(N8779) );
  CMX2X1 U24930 ( .A0(N8216), .A1(N8215), .S(n3875), .Z(n14140) );
  CMXI2X1 U24931 ( .A0(n14140), .A1(n14070), .S(n4171), .Z(n14207) );
  CMX2X1 U24932 ( .A0(n14071), .A1(n14207), .S(n4371), .Z(n14340) );
  CMXI2X1 U24933 ( .A0(n14072), .A1(n14340), .S(n3350), .Z(N8329) );
  CMXI2X1 U24934 ( .A0(n4424), .A1(n14074), .S(n3780), .Z(n14076) );
  CMXI2X1 U24935 ( .A0(n14076), .A1(n14075), .S(n3350), .Z(N8284) );
  CMX2X1 U24936 ( .A0(N7765), .A1(N7764), .S(n3876), .Z(n14083) );
  CMXI2X1 U24937 ( .A0(n14083), .A1(n14077), .S(n4171), .Z(n14090) );
  CMX2X1 U24938 ( .A0(n14078), .A1(n14090), .S(n4330), .Z(n14103) );
  CMXI2X1 U24939 ( .A0(n14079), .A1(n14103), .S(n3350), .Z(N8780) );
  CMX2X1 U24940 ( .A0(N7764), .A1(N7763), .S(n3877), .Z(n14086) );
  CMXI2X1 U24941 ( .A0(n14086), .A1(n14080), .S(n4171), .Z(n14093) );
  CMX2X1 U24942 ( .A0(n14081), .A1(n14093), .S(n4369), .Z(n14106) );
  CMXI2X1 U24943 ( .A0(n14082), .A1(n14106), .S(n3350), .Z(N8781) );
  CMX2X1 U24944 ( .A0(N7763), .A1(N7762), .S(n3878), .Z(n14089) );
  CMXI2X1 U24945 ( .A0(n14089), .A1(n14083), .S(n4170), .Z(n14096) );
  CMX2X1 U24946 ( .A0(n14084), .A1(n14096), .S(n4373), .Z(n14112) );
  CMXI2X1 U24947 ( .A0(n14085), .A1(n14112), .S(n3350), .Z(N8782) );
  CMX2X1 U24948 ( .A0(N7762), .A1(N7761), .S(n3879), .Z(n14092) );
  CMXI2X1 U24949 ( .A0(n14092), .A1(n14086), .S(n4170), .Z(n14099) );
  CMX2X1 U24950 ( .A0(n14087), .A1(n14099), .S(n4372), .Z(n14115) );
  CMXI2X1 U24951 ( .A0(n14088), .A1(n14115), .S(n3350), .Z(N8783) );
  CMX2X1 U24952 ( .A0(N7761), .A1(N7760), .S(n3880), .Z(n14095) );
  CMXI2X1 U24953 ( .A0(n14095), .A1(n14089), .S(n4170), .Z(n14102) );
  CMX2X1 U24954 ( .A0(n14090), .A1(n14102), .S(n4368), .Z(n14118) );
  CMXI2X1 U24955 ( .A0(n14091), .A1(n14118), .S(n3353), .Z(N8784) );
  CMX2X1 U24956 ( .A0(N7760), .A1(N7759), .S(n3870), .Z(n14098) );
  CMXI2X1 U24957 ( .A0(n14098), .A1(n14092), .S(n4170), .Z(n14105) );
  CMX2X1 U24958 ( .A0(n14093), .A1(n14105), .S(n4374), .Z(n14121) );
  CMXI2X1 U24959 ( .A0(n14094), .A1(n14121), .S(n3353), .Z(N8785) );
  CMX2X1 U24960 ( .A0(N7759), .A1(N7758), .S(n3871), .Z(n14101) );
  CMXI2X1 U24961 ( .A0(n14101), .A1(n14095), .S(n4170), .Z(n14111) );
  CMX2X1 U24962 ( .A0(n14096), .A1(n14111), .S(n4375), .Z(n14124) );
  CMXI2X1 U24963 ( .A0(n14097), .A1(n14124), .S(n3353), .Z(N8786) );
  CMX2X1 U24964 ( .A0(N7758), .A1(N7757), .S(n3872), .Z(n14104) );
  CMXI2X1 U24965 ( .A0(n14104), .A1(n14098), .S(n4170), .Z(n14114) );
  CMX2X1 U24966 ( .A0(n14099), .A1(n14114), .S(n4365), .Z(n14127) );
  CMXI2X1 U24967 ( .A0(n14100), .A1(n14127), .S(n3353), .Z(N8787) );
  CMX2X1 U24968 ( .A0(N7757), .A1(N7756), .S(n3873), .Z(n14110) );
  CMXI2X1 U24969 ( .A0(n14110), .A1(n14101), .S(n4170), .Z(n14117) );
  CMX2X1 U24970 ( .A0(n14102), .A1(n14117), .S(n4366), .Z(n14130) );
  CMXI2X1 U24971 ( .A0(n14103), .A1(n14130), .S(n3353), .Z(N8788) );
  CMX2X1 U24972 ( .A0(N7756), .A1(N7755), .S(n3863), .Z(n14113) );
  CMXI2X1 U24973 ( .A0(n14113), .A1(n14104), .S(n4170), .Z(n14120) );
  CMX2X1 U24974 ( .A0(n14105), .A1(n14120), .S(n4370), .Z(n14133) );
  CMXI2X1 U24975 ( .A0(n14106), .A1(n14133), .S(n3353), .Z(N8789) );
  CMX2X1 U24976 ( .A0(N8215), .A1(N8214), .S(n3877), .Z(n14173) );
  CMXI2X1 U24977 ( .A0(n14173), .A1(n14107), .S(n4170), .Z(n14240) );
  CMX2X1 U24978 ( .A0(n14108), .A1(n14240), .S(n4366), .Z(n14373) );
  CMXI2X1 U24979 ( .A0(n14109), .A1(n14373), .S(n3353), .Z(N8330) );
  CMX2X1 U24980 ( .A0(N7755), .A1(N7754), .S(n3878), .Z(n14116) );
  CMXI2X1 U24981 ( .A0(n14116), .A1(n14110), .S(n4170), .Z(n14123) );
  CMX2X1 U24982 ( .A0(n14111), .A1(n14123), .S(n4370), .Z(n14136) );
  CMXI2X1 U24983 ( .A0(n14112), .A1(n14136), .S(n3352), .Z(N8790) );
  CMX2X1 U24984 ( .A0(N7754), .A1(N7753), .S(n3879), .Z(n14119) );
  CMXI2X1 U24985 ( .A0(n14119), .A1(n14113), .S(n4170), .Z(n14126) );
  CMX2X1 U24986 ( .A0(n14114), .A1(n14126), .S(n4367), .Z(n14139) );
  CMXI2X1 U24987 ( .A0(n14115), .A1(n14139), .S(n3352), .Z(N8791) );
  CMX2X1 U24988 ( .A0(N7753), .A1(N7752), .S(n3880), .Z(n14122) );
  CMXI2X1 U24989 ( .A0(n14122), .A1(n14116), .S(n4170), .Z(n14129) );
  CMX2X1 U24990 ( .A0(n14117), .A1(n14129), .S(n4339), .Z(n14145) );
  CMXI2X1 U24991 ( .A0(n14118), .A1(n14145), .S(n3352), .Z(N8792) );
  CMX2X1 U24992 ( .A0(N7752), .A1(N7751), .S(n3881), .Z(n14125) );
  CMXI2X1 U24993 ( .A0(n14125), .A1(n14119), .S(n4170), .Z(n14132) );
  CMX2X1 U24994 ( .A0(n14120), .A1(n14132), .S(n4340), .Z(n14148) );
  CMXI2X1 U24995 ( .A0(n14121), .A1(n14148), .S(n3352), .Z(N8793) );
  CMX2X1 U24996 ( .A0(N7751), .A1(N7750), .S(n3862), .Z(n14128) );
  CMXI2X1 U24997 ( .A0(n14128), .A1(n14122), .S(n4170), .Z(n14135) );
  CMX2X1 U24998 ( .A0(n14123), .A1(n14135), .S(n4331), .Z(n14151) );
  CMXI2X1 U24999 ( .A0(n14124), .A1(n14151), .S(n3352), .Z(N8794) );
  CMX2X1 U25000 ( .A0(N7750), .A1(N7749), .S(n3863), .Z(n14131) );
  CMXI2X1 U25001 ( .A0(n14131), .A1(n14125), .S(n4170), .Z(n14138) );
  CMX2X1 U25002 ( .A0(n14126), .A1(n14138), .S(n4332), .Z(n14154) );
  CMXI2X1 U25003 ( .A0(n14127), .A1(n14154), .S(n3352), .Z(N8795) );
  CMX2X1 U25004 ( .A0(N7749), .A1(N7748), .S(n3865), .Z(n14134) );
  CMXI2X1 U25005 ( .A0(n14134), .A1(n14128), .S(n4170), .Z(n14144) );
  CMX2X1 U25006 ( .A0(n14129), .A1(n14144), .S(n4333), .Z(n14157) );
  CMXI2X1 U25007 ( .A0(n14130), .A1(n14157), .S(n3352), .Z(N8796) );
  CMX2X1 U25008 ( .A0(N7748), .A1(N7747), .S(n3866), .Z(n14137) );
  CMXI2X1 U25009 ( .A0(n14137), .A1(n14131), .S(n4169), .Z(n14147) );
  CMX2X1 U25010 ( .A0(n14132), .A1(n14147), .S(n4336), .Z(n14160) );
  CMXI2X1 U25011 ( .A0(n14133), .A1(n14160), .S(n3352), .Z(N8797) );
  CMX2X1 U25012 ( .A0(N7747), .A1(N7746), .S(n3864), .Z(n14143) );
  CMXI2X1 U25013 ( .A0(n14143), .A1(n14134), .S(n4169), .Z(n14150) );
  CMX2X1 U25014 ( .A0(n14135), .A1(n14150), .S(n4337), .Z(n14163) );
  CMXI2X1 U25015 ( .A0(n14136), .A1(n14163), .S(n3352), .Z(N8798) );
  CMX2X1 U25016 ( .A0(N7746), .A1(N7745), .S(n3865), .Z(n14146) );
  CMXI2X1 U25017 ( .A0(n14146), .A1(n14137), .S(n4169), .Z(n14153) );
  CMX2X1 U25018 ( .A0(n14138), .A1(n14153), .S(n4338), .Z(n14166) );
  CMXI2X1 U25019 ( .A0(n14139), .A1(n14166), .S(n3352), .Z(N8799) );
  CMX2X1 U25020 ( .A0(N8214), .A1(N8213), .S(n3881), .Z(n14206) );
  CMXI2X1 U25021 ( .A0(n14206), .A1(n14140), .S(n4169), .Z(n14273) );
  CMX2X1 U25022 ( .A0(n14141), .A1(n14273), .S(n4371), .Z(n14406) );
  CMXI2X1 U25023 ( .A0(n14142), .A1(n14406), .S(n3352), .Z(N8331) );
  CMX2X1 U25024 ( .A0(N7745), .A1(N7744), .S(n3862), .Z(n14149) );
  CMXI2X1 U25025 ( .A0(n14149), .A1(n14143), .S(n4169), .Z(n14156) );
  CMX2X1 U25026 ( .A0(n14144), .A1(n14156), .S(n4366), .Z(n14169) );
  CMXI2X1 U25027 ( .A0(n14145), .A1(n14169), .S(n3355), .Z(N8800) );
  CMX2X1 U25028 ( .A0(N7744), .A1(N7743), .S(n3863), .Z(n14152) );
  CMXI2X1 U25029 ( .A0(n14152), .A1(n14146), .S(n4169), .Z(n14159) );
  CMX2X1 U25030 ( .A0(n14147), .A1(n14159), .S(n4370), .Z(n14172) );
  CMXI2X1 U25031 ( .A0(n14148), .A1(n14172), .S(n3355), .Z(N8801) );
  CMX2X1 U25032 ( .A0(N7743), .A1(N7742), .S(n3878), .Z(n14155) );
  CMXI2X1 U25033 ( .A0(n14155), .A1(n14149), .S(n4169), .Z(n14162) );
  CMX2X1 U25034 ( .A0(n14150), .A1(n14162), .S(n4372), .Z(n14178) );
  CMXI2X1 U25035 ( .A0(n14151), .A1(n14178), .S(n3355), .Z(N8802) );
  CMX2X1 U25036 ( .A0(N7742), .A1(N7741), .S(n3876), .Z(n14158) );
  CMXI2X1 U25037 ( .A0(n14158), .A1(n14152), .S(n4169), .Z(n14165) );
  CMX2X1 U25038 ( .A0(n14153), .A1(n14165), .S(n4368), .Z(n14181) );
  CMXI2X1 U25039 ( .A0(n14154), .A1(n14181), .S(n3354), .Z(N8803) );
  CMX2X1 U25040 ( .A0(N7741), .A1(N7740), .S(n3877), .Z(n14161) );
  CMXI2X1 U25041 ( .A0(n14161), .A1(n14155), .S(n4169), .Z(n14168) );
  CMX2X1 U25042 ( .A0(n14156), .A1(n14168), .S(n4375), .Z(n14184) );
  CMXI2X1 U25043 ( .A0(n14157), .A1(n14184), .S(n3354), .Z(N8804) );
  CMX2X1 U25044 ( .A0(N7740), .A1(N7739), .S(n3879), .Z(n14164) );
  CMXI2X1 U25045 ( .A0(n14164), .A1(n14158), .S(n4169), .Z(n14171) );
  CMX2X1 U25046 ( .A0(n14159), .A1(n14171), .S(n4365), .Z(n14187) );
  CMXI2X1 U25047 ( .A0(n14160), .A1(n14187), .S(n3354), .Z(N8805) );
  CMX2X1 U25048 ( .A0(N7739), .A1(N7738), .S(n3880), .Z(n14167) );
  CMXI2X1 U25049 ( .A0(n14167), .A1(n14161), .S(n4169), .Z(n14177) );
  CMX2X1 U25050 ( .A0(n14162), .A1(n14177), .S(n4369), .Z(n14190) );
  CMXI2X1 U25051 ( .A0(n14163), .A1(n14190), .S(n3354), .Z(N8806) );
  CMX2X1 U25052 ( .A0(N7738), .A1(N7737), .S(n3877), .Z(n14170) );
  CMXI2X1 U25053 ( .A0(n14170), .A1(n14164), .S(n4169), .Z(n14180) );
  CMX2X1 U25054 ( .A0(n14165), .A1(n14180), .S(n4374), .Z(n14193) );
  CMXI2X1 U25055 ( .A0(n14166), .A1(n14193), .S(n3354), .Z(N8807) );
  CMX2X1 U25056 ( .A0(N7737), .A1(N7736), .S(n3878), .Z(n14176) );
  CMXI2X1 U25057 ( .A0(n14176), .A1(n14167), .S(n4169), .Z(n14183) );
  CMX2X1 U25058 ( .A0(n14168), .A1(n14183), .S(n4373), .Z(n14196) );
  CMXI2X1 U25059 ( .A0(n14169), .A1(n14196), .S(n3354), .Z(N8808) );
  CMX2X1 U25060 ( .A0(N7736), .A1(N7735), .S(n3879), .Z(n14179) );
  CMXI2X1 U25061 ( .A0(n14179), .A1(n14170), .S(n4169), .Z(n14186) );
  CMX2X1 U25062 ( .A0(n14171), .A1(n14186), .S(n4371), .Z(n14199) );
  CMXI2X1 U25063 ( .A0(n14172), .A1(n14199), .S(n3354), .Z(N8809) );
  CMX2X1 U25064 ( .A0(N8213), .A1(N8212), .S(n3880), .Z(n14239) );
  CMXI2X1 U25065 ( .A0(n14239), .A1(n14173), .S(n4169), .Z(n14306) );
  CMX2X1 U25066 ( .A0(n14174), .A1(n14306), .S(n4318), .Z(n14443) );
  CMXI2X1 U25067 ( .A0(n14175), .A1(n14443), .S(n3354), .Z(N8332) );
  CMX2X1 U25068 ( .A0(N7735), .A1(N7734), .S(n3875), .Z(n14182) );
  CMXI2X1 U25069 ( .A0(n14182), .A1(n14176), .S(n4169), .Z(n14189) );
  CMX2X1 U25070 ( .A0(n14177), .A1(n14189), .S(n4318), .Z(n14202) );
  CMXI2X1 U25071 ( .A0(n14178), .A1(n14202), .S(n3354), .Z(N8810) );
  CMX2X1 U25072 ( .A0(N7734), .A1(N7733), .S(n3876), .Z(n14185) );
  CMXI2X1 U25073 ( .A0(n14185), .A1(n14179), .S(n4168), .Z(n14192) );
  CMX2X1 U25074 ( .A0(n14180), .A1(n14192), .S(n4318), .Z(n14205) );
  CMXI2X1 U25075 ( .A0(n14181), .A1(n14205), .S(n3354), .Z(N8811) );
  CMX2X1 U25076 ( .A0(N7733), .A1(N7732), .S(n3877), .Z(n14188) );
  CMXI2X1 U25077 ( .A0(n14188), .A1(n14182), .S(n4168), .Z(n14195) );
  CMX2X1 U25078 ( .A0(n14183), .A1(n14195), .S(n4318), .Z(n14211) );
  CMXI2X1 U25079 ( .A0(n14184), .A1(n14211), .S(n3354), .Z(N8812) );
  CMX2X1 U25080 ( .A0(N7732), .A1(N7731), .S(n3878), .Z(n14191) );
  CMXI2X1 U25081 ( .A0(n14191), .A1(n14185), .S(n4168), .Z(n14198) );
  CMX2X1 U25082 ( .A0(n14186), .A1(n14198), .S(n4318), .Z(n14214) );
  CMXI2X1 U25083 ( .A0(n14187), .A1(n14214), .S(n3353), .Z(N8813) );
  CMX2X1 U25084 ( .A0(N7731), .A1(N7730), .S(n3865), .Z(n14194) );
  CMXI2X1 U25085 ( .A0(n14194), .A1(n14188), .S(n4168), .Z(n14201) );
  CMX2X1 U25086 ( .A0(n14189), .A1(n14201), .S(n4318), .Z(n14217) );
  CMXI2X1 U25087 ( .A0(n14190), .A1(n14217), .S(n3353), .Z(N8814) );
  CMX2X1 U25088 ( .A0(N7730), .A1(N7729), .S(n3881), .Z(n14197) );
  CMXI2X1 U25089 ( .A0(n14197), .A1(n14191), .S(n4168), .Z(n14204) );
  CMX2X1 U25090 ( .A0(n14192), .A1(n14204), .S(n4318), .Z(n14220) );
  CMXI2X1 U25091 ( .A0(n14193), .A1(n14220), .S(n3353), .Z(N8815) );
  CMX2X1 U25092 ( .A0(N7729), .A1(N7728), .S(n3862), .Z(n14200) );
  CMXI2X1 U25093 ( .A0(n14200), .A1(n14194), .S(n4168), .Z(n14210) );
  CMX2X1 U25094 ( .A0(n14195), .A1(n14210), .S(n4318), .Z(n14223) );
  CMXI2X1 U25095 ( .A0(n14196), .A1(n14223), .S(n3353), .Z(N8816) );
  CMX2X1 U25096 ( .A0(N7728), .A1(N7727), .S(n3863), .Z(n14203) );
  CMXI2X1 U25097 ( .A0(n14203), .A1(n14197), .S(n4168), .Z(n14213) );
  CMX2X1 U25098 ( .A0(n14198), .A1(n14213), .S(n4318), .Z(n14226) );
  CMXI2X1 U25099 ( .A0(n14199), .A1(n14226), .S(n3356), .Z(N8817) );
  CMX2X1 U25100 ( .A0(N7727), .A1(N7726), .S(n3864), .Z(n14209) );
  CMXI2X1 U25101 ( .A0(n14209), .A1(n14200), .S(n4168), .Z(n14216) );
  CMX2X1 U25102 ( .A0(n14201), .A1(n14216), .S(n4318), .Z(n14229) );
  CMXI2X1 U25103 ( .A0(n14202), .A1(n14229), .S(n3356), .Z(N8818) );
  CMX2X1 U25104 ( .A0(N7726), .A1(N7725), .S(n3865), .Z(n14212) );
  CMXI2X1 U25105 ( .A0(n14212), .A1(n14203), .S(n4168), .Z(n14219) );
  CMX2X1 U25106 ( .A0(n14204), .A1(n14219), .S(n4318), .Z(n14232) );
  CMXI2X1 U25107 ( .A0(n14205), .A1(n14232), .S(n3356), .Z(N8819) );
  CMX2X1 U25108 ( .A0(N8212), .A1(N8211), .S(n3866), .Z(n14272) );
  CMXI2X1 U25109 ( .A0(n14272), .A1(n14206), .S(n4168), .Z(n14339) );
  CMX2X1 U25110 ( .A0(n14207), .A1(n14339), .S(n4317), .Z(n14476) );
  CMXI2X1 U25111 ( .A0(n14208), .A1(n14476), .S(n3356), .Z(N8333) );
  CMX2X1 U25112 ( .A0(N7725), .A1(N7724), .S(n3867), .Z(n14215) );
  CMXI2X1 U25113 ( .A0(n14215), .A1(n14209), .S(n4168), .Z(n14222) );
  CMX2X1 U25114 ( .A0(n14210), .A1(n14222), .S(n4317), .Z(n14235) );
  CMXI2X1 U25115 ( .A0(n14211), .A1(n14235), .S(n3356), .Z(N8820) );
  CMX2X1 U25116 ( .A0(N7724), .A1(N7723), .S(n3879), .Z(n14218) );
  CMXI2X1 U25117 ( .A0(n14218), .A1(n14212), .S(n4168), .Z(n14225) );
  CMX2X1 U25118 ( .A0(n14213), .A1(n14225), .S(n4317), .Z(n14238) );
  CMXI2X1 U25119 ( .A0(n14214), .A1(n14238), .S(n3356), .Z(N8821) );
  CMX2X1 U25120 ( .A0(N7723), .A1(N7722), .S(n3868), .Z(n14221) );
  CMXI2X1 U25121 ( .A0(n14221), .A1(n14215), .S(n4168), .Z(n14228) );
  CMX2X1 U25122 ( .A0(n14216), .A1(n14228), .S(n4317), .Z(n14244) );
  CMXI2X1 U25123 ( .A0(n14217), .A1(n14244), .S(n3356), .Z(N8822) );
  CMX2X1 U25124 ( .A0(N7722), .A1(N7721), .S(n3869), .Z(n14224) );
  CMXI2X1 U25125 ( .A0(n14224), .A1(n14218), .S(n4168), .Z(n14231) );
  CMX2X1 U25126 ( .A0(n14219), .A1(n14231), .S(n4317), .Z(n14247) );
  CMXI2X1 U25127 ( .A0(n14220), .A1(n14247), .S(n3356), .Z(N8823) );
  CMX2X1 U25128 ( .A0(N7721), .A1(N7720), .S(n3881), .Z(n14227) );
  CMXI2X1 U25129 ( .A0(n14227), .A1(n14221), .S(n4168), .Z(n14234) );
  CMX2X1 U25130 ( .A0(n14222), .A1(n14234), .S(n4317), .Z(n14250) );
  CMXI2X1 U25131 ( .A0(n14223), .A1(n14250), .S(n3356), .Z(N8824) );
  CMX2X1 U25132 ( .A0(N7720), .A1(N7719), .S(n3862), .Z(n14230) );
  CMXI2X1 U25133 ( .A0(n14230), .A1(n14224), .S(n4168), .Z(n14237) );
  CMX2X1 U25134 ( .A0(n14225), .A1(n14237), .S(n4317), .Z(n14253) );
  CMXI2X1 U25135 ( .A0(n14226), .A1(n14253), .S(n3356), .Z(N8825) );
  CMX2X1 U25136 ( .A0(N7719), .A1(N7718), .S(n3863), .Z(n14233) );
  CMXI2X1 U25137 ( .A0(n14233), .A1(n14227), .S(n4167), .Z(n14243) );
  CMX2X1 U25138 ( .A0(n14228), .A1(n14243), .S(n4317), .Z(n14256) );
  CMXI2X1 U25139 ( .A0(n14229), .A1(n14256), .S(n3355), .Z(N8826) );
  CMX2X1 U25140 ( .A0(N7718), .A1(N7717), .S(n3864), .Z(n14236) );
  CMXI2X1 U25141 ( .A0(n14236), .A1(n14230), .S(n4167), .Z(n14246) );
  CMX2X1 U25142 ( .A0(n14231), .A1(n14246), .S(n4317), .Z(n14259) );
  CMXI2X1 U25143 ( .A0(n14232), .A1(n14259), .S(n3355), .Z(N8827) );
  CMX2X1 U25144 ( .A0(N7717), .A1(N7716), .S(n3879), .Z(n14242) );
  CMXI2X1 U25145 ( .A0(n14242), .A1(n14233), .S(n4167), .Z(n14249) );
  CMX2X1 U25146 ( .A0(n14234), .A1(n14249), .S(n4317), .Z(n14262) );
  CMXI2X1 U25147 ( .A0(n14235), .A1(n14262), .S(n3355), .Z(N8828) );
  CMX2X1 U25148 ( .A0(N7716), .A1(N7715), .S(n3880), .Z(n14245) );
  CMXI2X1 U25149 ( .A0(n14245), .A1(n14236), .S(n4167), .Z(n14252) );
  CMX2X1 U25150 ( .A0(n14237), .A1(n14252), .S(n4317), .Z(n14265) );
  CMXI2X1 U25151 ( .A0(n14238), .A1(n14265), .S(n3355), .Z(N8829) );
  CMX2X1 U25152 ( .A0(N8211), .A1(N8210), .S(n3881), .Z(n14305) );
  CMXI2X1 U25153 ( .A0(n14305), .A1(n14239), .S(n4167), .Z(n14372) );
  CMX2X1 U25154 ( .A0(n14240), .A1(n14372), .S(n4316), .Z(n14509) );
  CMXI2X1 U25155 ( .A0(n14241), .A1(n14509), .S(n3355), .Z(N8334) );
  CMX2X1 U25156 ( .A0(N7715), .A1(N7714), .S(n3862), .Z(n14248) );
  CMXI2X1 U25157 ( .A0(n14248), .A1(n14242), .S(n4167), .Z(n14255) );
  CMX2X1 U25158 ( .A0(n14243), .A1(n14255), .S(n4316), .Z(n14268) );
  CMXI2X1 U25159 ( .A0(n14244), .A1(n14268), .S(n3355), .Z(N8830) );
  CMX2X1 U25160 ( .A0(N7714), .A1(N7713), .S(n3866), .Z(n14251) );
  CMXI2X1 U25161 ( .A0(n14251), .A1(n14245), .S(n4167), .Z(n14258) );
  CMX2X1 U25162 ( .A0(n14246), .A1(n14258), .S(n4316), .Z(n14271) );
  CMXI2X1 U25163 ( .A0(n14247), .A1(n14271), .S(n3355), .Z(N8831) );
  CMX2X1 U25164 ( .A0(N7713), .A1(N7712), .S(n3870), .Z(n14254) );
  CMXI2X1 U25165 ( .A0(n14254), .A1(n14248), .S(n4167), .Z(n14261) );
  CMX2X1 U25166 ( .A0(n14249), .A1(n14261), .S(n4316), .Z(n14277) );
  CMXI2X1 U25167 ( .A0(n14250), .A1(n14277), .S(n3355), .Z(N8832) );
  CMX2X1 U25168 ( .A0(N7712), .A1(N7711), .S(n3871), .Z(n14257) );
  CMXI2X1 U25169 ( .A0(n14257), .A1(n14251), .S(n4167), .Z(n14264) );
  CMX2X1 U25170 ( .A0(n14252), .A1(n14264), .S(n4316), .Z(n14280) );
  CMXI2X1 U25171 ( .A0(n14253), .A1(n14280), .S(n3358), .Z(N8833) );
  CMX2X1 U25172 ( .A0(N7711), .A1(N7710), .S(n3872), .Z(n14260) );
  CMXI2X1 U25173 ( .A0(n14260), .A1(n14254), .S(n4167), .Z(n14267) );
  CMX2X1 U25174 ( .A0(n14255), .A1(n14267), .S(n4316), .Z(n14283) );
  CMXI2X1 U25175 ( .A0(n14256), .A1(n14283), .S(n3358), .Z(N8834) );
  CMX2X1 U25176 ( .A0(N7710), .A1(N7709), .S(n3873), .Z(n14263) );
  CMXI2X1 U25177 ( .A0(n14263), .A1(n14257), .S(n4167), .Z(n14270) );
  CMX2X1 U25178 ( .A0(n14258), .A1(n14270), .S(n4316), .Z(n14286) );
  CMXI2X1 U25179 ( .A0(n14259), .A1(n14286), .S(n3358), .Z(N8835) );
  CMX2X1 U25180 ( .A0(N7709), .A1(N7708), .S(n3874), .Z(n14266) );
  CMXI2X1 U25181 ( .A0(n14266), .A1(n14260), .S(n4167), .Z(n14276) );
  CMX2X1 U25182 ( .A0(n14261), .A1(n14276), .S(n4316), .Z(n14289) );
  CMXI2X1 U25183 ( .A0(n14262), .A1(n14289), .S(n3358), .Z(N8836) );
  CMX2X1 U25184 ( .A0(N7708), .A1(N7707), .S(n3875), .Z(n14269) );
  CMXI2X1 U25185 ( .A0(n14269), .A1(n14263), .S(n4167), .Z(n14279) );
  CMX2X1 U25186 ( .A0(n14264), .A1(n14279), .S(n4316), .Z(n14292) );
  CMXI2X1 U25187 ( .A0(n14265), .A1(n14292), .S(n3358), .Z(N8837) );
  CMX2X1 U25188 ( .A0(N7707), .A1(N7706), .S(n3876), .Z(n14275) );
  CMXI2X1 U25189 ( .A0(n14275), .A1(n14266), .S(n4167), .Z(n14282) );
  CMX2X1 U25190 ( .A0(n14267), .A1(n14282), .S(n4316), .Z(n14295) );
  CMXI2X1 U25191 ( .A0(n14268), .A1(n14295), .S(n3358), .Z(N8838) );
  CMX2X1 U25192 ( .A0(N7706), .A1(N7705), .S(n3880), .Z(n14278) );
  CMXI2X1 U25193 ( .A0(n14278), .A1(n14269), .S(n4167), .Z(n14285) );
  CMX2X1 U25194 ( .A0(n14270), .A1(n14285), .S(n4315), .Z(n14298) );
  CMXI2X1 U25195 ( .A0(n14271), .A1(n14298), .S(n3358), .Z(N8839) );
  CMX2X1 U25196 ( .A0(N8210), .A1(N8209), .S(n3881), .Z(n14338) );
  CMXI2X1 U25197 ( .A0(n14338), .A1(n14272), .S(n4167), .Z(n14405) );
  CMX2X1 U25198 ( .A0(n14273), .A1(n14405), .S(n4315), .Z(n14542) );
  CMXI2X1 U25199 ( .A0(n14274), .A1(n14542), .S(n3357), .Z(N8335) );
  CMX2X1 U25200 ( .A0(N7705), .A1(N7704), .S(n3877), .Z(n14281) );
  CMXI2X1 U25201 ( .A0(n14281), .A1(n14275), .S(n4166), .Z(n14288) );
  CMX2X1 U25202 ( .A0(n14276), .A1(n14288), .S(n4315), .Z(n14301) );
  CMXI2X1 U25203 ( .A0(n14277), .A1(n14301), .S(n3357), .Z(N8840) );
  CMX2X1 U25204 ( .A0(N7704), .A1(N7703), .S(n3878), .Z(n14284) );
  CMXI2X1 U25205 ( .A0(n14284), .A1(n14278), .S(n4166), .Z(n14291) );
  CMX2X1 U25206 ( .A0(n14279), .A1(n14291), .S(n4315), .Z(n14304) );
  CMXI2X1 U25207 ( .A0(n14280), .A1(n14304), .S(n3357), .Z(N8841) );
  CMX2X1 U25208 ( .A0(N7703), .A1(N7702), .S(n3865), .Z(n14287) );
  CMXI2X1 U25209 ( .A0(n14287), .A1(n14281), .S(n4166), .Z(n14294) );
  CMX2X1 U25210 ( .A0(n14282), .A1(n14294), .S(n4315), .Z(n14310) );
  CMXI2X1 U25211 ( .A0(n14283), .A1(n14310), .S(n3357), .Z(N8842) );
  CMX2X1 U25212 ( .A0(N7702), .A1(N7701), .S(n3866), .Z(n14290) );
  CMXI2X1 U25213 ( .A0(n14290), .A1(n14284), .S(n4166), .Z(n14297) );
  CMX2X1 U25214 ( .A0(n14285), .A1(n14297), .S(n4315), .Z(n14313) );
  CMXI2X1 U25215 ( .A0(n14286), .A1(n14313), .S(n3357), .Z(N8843) );
  CMX2X1 U25216 ( .A0(N7701), .A1(N7700), .S(n3867), .Z(n14293) );
  CMXI2X1 U25217 ( .A0(n14293), .A1(n14287), .S(n4166), .Z(n14300) );
  CMX2X1 U25218 ( .A0(n14288), .A1(n14300), .S(n4315), .Z(n14316) );
  CMXI2X1 U25219 ( .A0(n14289), .A1(n14316), .S(n3357), .Z(N8844) );
  CMX2X1 U25220 ( .A0(N7700), .A1(N7699), .S(n3868), .Z(n14296) );
  CMXI2X1 U25221 ( .A0(n14296), .A1(n14290), .S(n4166), .Z(n14303) );
  CMX2X1 U25222 ( .A0(n14291), .A1(n14303), .S(n4315), .Z(n14319) );
  CMXI2X1 U25223 ( .A0(n14292), .A1(n14319), .S(n3357), .Z(N8845) );
  CMX2X1 U25224 ( .A0(N7699), .A1(N7698), .S(n3863), .Z(n14299) );
  CMXI2X1 U25225 ( .A0(n14299), .A1(n14293), .S(n4166), .Z(n14309) );
  CMX2X1 U25226 ( .A0(n14294), .A1(n14309), .S(n4315), .Z(n14322) );
  CMXI2X1 U25227 ( .A0(n14295), .A1(n14322), .S(n3357), .Z(N8846) );
  CMX2X1 U25228 ( .A0(N7698), .A1(N7697), .S(n3864), .Z(n14302) );
  CMXI2X1 U25229 ( .A0(n14302), .A1(n14296), .S(n4166), .Z(n14312) );
  CMX2X1 U25230 ( .A0(n14297), .A1(n14312), .S(n4315), .Z(n14325) );
  CMXI2X1 U25231 ( .A0(n14298), .A1(n14325), .S(n3357), .Z(N8847) );
  CMX2X1 U25232 ( .A0(N7697), .A1(N7696), .S(n3865), .Z(n14308) );
  CMXI2X1 U25233 ( .A0(n14308), .A1(n14299), .S(n4166), .Z(n14315) );
  CMX2X1 U25234 ( .A0(n14300), .A1(n14315), .S(n4315), .Z(n14328) );
  CMXI2X1 U25235 ( .A0(n14301), .A1(n14328), .S(n3357), .Z(N8848) );
  CMX2X1 U25236 ( .A0(N7696), .A1(N7695), .S(n3866), .Z(n14311) );
  CMXI2X1 U25237 ( .A0(n14311), .A1(n14302), .S(n4166), .Z(n14318) );
  CMX2X1 U25238 ( .A0(n14303), .A1(n14318), .S(n4314), .Z(n14331) );
  CMXI2X1 U25239 ( .A0(n14304), .A1(n14331), .S(n3360), .Z(N8849) );
  CMX2X1 U25240 ( .A0(N8209), .A1(N8208), .S(n3867), .Z(n14371) );
  CMXI2X1 U25241 ( .A0(n14371), .A1(n14305), .S(n4166), .Z(n14442) );
  CMX2X1 U25242 ( .A0(n14306), .A1(n14442), .S(n4314), .Z(n14575) );
  CMXI2X1 U25243 ( .A0(n14307), .A1(n14575), .S(n3360), .Z(N8336) );
  CMX2X1 U25244 ( .A0(N7695), .A1(N7694), .S(n3879), .Z(n14314) );
  CMXI2X1 U25245 ( .A0(n14314), .A1(n14308), .S(n4166), .Z(n14321) );
  CMX2X1 U25246 ( .A0(n14309), .A1(n14321), .S(n4314), .Z(n14334) );
  CMXI2X1 U25247 ( .A0(n14310), .A1(n14334), .S(n3360), .Z(N8850) );
  CMX2X1 U25248 ( .A0(N7694), .A1(N7693), .S(n3880), .Z(n14317) );
  CMXI2X1 U25249 ( .A0(n14317), .A1(n14311), .S(n4166), .Z(n14324) );
  CMX2X1 U25250 ( .A0(n14312), .A1(n14324), .S(n4314), .Z(n14337) );
  CMXI2X1 U25251 ( .A0(n14313), .A1(n14337), .S(n3359), .Z(N8851) );
  CMX2X1 U25252 ( .A0(N7693), .A1(N7692), .S(n3881), .Z(n14320) );
  CMXI2X1 U25253 ( .A0(n14320), .A1(n14314), .S(n4166), .Z(n14327) );
  CMX2X1 U25254 ( .A0(n14315), .A1(n14327), .S(n4314), .Z(n14343) );
  CMXI2X1 U25255 ( .A0(n14316), .A1(n14343), .S(n3359), .Z(N8852) );
  CMX2X1 U25256 ( .A0(N7692), .A1(N7691), .S(n3862), .Z(n14323) );
  CMXI2X1 U25257 ( .A0(n14323), .A1(n14317), .S(n4166), .Z(n14330) );
  CMX2X1 U25258 ( .A0(n14318), .A1(n14330), .S(n4314), .Z(n14346) );
  CMXI2X1 U25259 ( .A0(n14319), .A1(n14346), .S(n3359), .Z(N8853) );
  CMX2X1 U25260 ( .A0(N7691), .A1(N7690), .S(n3863), .Z(n14326) );
  CMXI2X1 U25261 ( .A0(n14326), .A1(n14320), .S(n4166), .Z(n14333) );
  CMX2X1 U25262 ( .A0(n14321), .A1(n14333), .S(n4314), .Z(n14349) );
  CMXI2X1 U25263 ( .A0(n14322), .A1(n14349), .S(n3359), .Z(N8854) );
  CMX2X1 U25264 ( .A0(N7690), .A1(N7689), .S(n3864), .Z(n14329) );
  CMXI2X1 U25265 ( .A0(n14329), .A1(n14323), .S(n4165), .Z(n14336) );
  CMX2X1 U25266 ( .A0(n14324), .A1(n14336), .S(n4314), .Z(n14352) );
  CMXI2X1 U25267 ( .A0(n14325), .A1(n14352), .S(n3359), .Z(N8855) );
  CMX2X1 U25268 ( .A0(N7689), .A1(N7688), .S(n3865), .Z(n14332) );
  CMXI2X1 U25269 ( .A0(n14332), .A1(n14326), .S(n4165), .Z(n14342) );
  CMX2X1 U25270 ( .A0(n14327), .A1(n14342), .S(n4314), .Z(n14355) );
  CMXI2X1 U25271 ( .A0(n14328), .A1(n14355), .S(n3359), .Z(N8856) );
  CMX2X1 U25272 ( .A0(N7688), .A1(N7687), .S(n3862), .Z(n14335) );
  CMXI2X1 U25273 ( .A0(n14335), .A1(n14329), .S(n4165), .Z(n14345) );
  CMX2X1 U25274 ( .A0(n14330), .A1(n14345), .S(n4314), .Z(n14358) );
  CMXI2X1 U25275 ( .A0(n14331), .A1(n14358), .S(n3359), .Z(N8857) );
  CMX2X1 U25276 ( .A0(N7687), .A1(N7686), .S(n3863), .Z(n14341) );
  CMXI2X1 U25277 ( .A0(n14341), .A1(n14332), .S(n4165), .Z(n14348) );
  CMX2X1 U25278 ( .A0(n14333), .A1(n14348), .S(n4314), .Z(n14361) );
  CMXI2X1 U25279 ( .A0(n14334), .A1(n14361), .S(n3359), .Z(N8858) );
  CMX2X1 U25280 ( .A0(N7686), .A1(N7685), .S(n3866), .Z(n14344) );
  CMXI2X1 U25281 ( .A0(n14344), .A1(n14335), .S(n4165), .Z(n14351) );
  CMX2X1 U25282 ( .A0(n14336), .A1(n14351), .S(n4313), .Z(n14364) );
  CMXI2X1 U25283 ( .A0(n14337), .A1(n14364), .S(n3359), .Z(N8859) );
  CMX2X1 U25284 ( .A0(N8208), .A1(N8207), .S(n3867), .Z(n14404) );
  CMXI2X1 U25285 ( .A0(n14404), .A1(n14338), .S(n4165), .Z(n14475) );
  CMX2X1 U25286 ( .A0(n14339), .A1(n14475), .S(n4313), .Z(n14608) );
  CMXI2X1 U25287 ( .A0(n14340), .A1(n14608), .S(n3359), .Z(N8337) );
  CMX2X1 U25288 ( .A0(N7685), .A1(N7684), .S(n3869), .Z(n14347) );
  CMXI2X1 U25289 ( .A0(n14347), .A1(n14341), .S(n4165), .Z(n14354) );
  CMX2X1 U25290 ( .A0(n14342), .A1(n14354), .S(n4313), .Z(n14367) );
  CMXI2X1 U25291 ( .A0(n14343), .A1(n14367), .S(n3359), .Z(N8860) );
  CMX2X1 U25292 ( .A0(N7684), .A1(N7683), .S(n3870), .Z(n14350) );
  CMXI2X1 U25293 ( .A0(n14350), .A1(n14344), .S(n4165), .Z(n14357) );
  CMX2X1 U25294 ( .A0(n14345), .A1(n14357), .S(n4313), .Z(n14370) );
  CMXI2X1 U25295 ( .A0(n14346), .A1(n14370), .S(n3358), .Z(N8861) );
  CMX2X1 U25296 ( .A0(N7683), .A1(N7682), .S(n3871), .Z(n14353) );
  CMXI2X1 U25297 ( .A0(n14353), .A1(n14347), .S(n4165), .Z(n14360) );
  CMX2X1 U25298 ( .A0(n14348), .A1(n14360), .S(n4313), .Z(n14376) );
  CMXI2X1 U25299 ( .A0(n14349), .A1(n14376), .S(n3358), .Z(N8862) );
  CMX2X1 U25300 ( .A0(N7682), .A1(N7681), .S(n3872), .Z(n14356) );
  CMXI2X1 U25301 ( .A0(n14356), .A1(n14350), .S(n4165), .Z(n14363) );
  CMX2X1 U25302 ( .A0(n14351), .A1(n14363), .S(n4313), .Z(n14379) );
  CMXI2X1 U25303 ( .A0(n14352), .A1(n14379), .S(n3358), .Z(N8863) );
  CMX2X1 U25304 ( .A0(N7681), .A1(N7680), .S(n3867), .Z(n14359) );
  CMXI2X1 U25305 ( .A0(n14359), .A1(n14353), .S(n4165), .Z(n14366) );
  CMX2X1 U25306 ( .A0(n14354), .A1(n14366), .S(n4313), .Z(n14382) );
  CMXI2X1 U25307 ( .A0(n14355), .A1(n14382), .S(n3358), .Z(N8864) );
  CMX2X1 U25308 ( .A0(N7680), .A1(N7679), .S(n3868), .Z(n14362) );
  CMXI2X1 U25309 ( .A0(n14362), .A1(n14356), .S(n4165), .Z(n14369) );
  CMX2X1 U25310 ( .A0(n14357), .A1(n14369), .S(n4313), .Z(n14385) );
  CMXI2X1 U25311 ( .A0(n14358), .A1(n14385), .S(n3361), .Z(N8865) );
  CMX2X1 U25312 ( .A0(N7679), .A1(N7678), .S(n3869), .Z(n14365) );
  CMXI2X1 U25313 ( .A0(n14365), .A1(n14359), .S(n4165), .Z(n14375) );
  CMX2X1 U25314 ( .A0(n14360), .A1(n14375), .S(n4313), .Z(n14388) );
  CMXI2X1 U25315 ( .A0(n14361), .A1(n14388), .S(n3361), .Z(N8866) );
  CMX2X1 U25316 ( .A0(N7678), .A1(N7677), .S(n3870), .Z(n14368) );
  CMXI2X1 U25317 ( .A0(n14368), .A1(n14362), .S(n4165), .Z(n14378) );
  CMX2X1 U25318 ( .A0(n14363), .A1(n14378), .S(n4313), .Z(n14391) );
  CMXI2X1 U25319 ( .A0(n14364), .A1(n14391), .S(n3361), .Z(N8867) );
  CMX2X1 U25320 ( .A0(N7677), .A1(N7676), .S(n3868), .Z(n14374) );
  CMXI2X1 U25321 ( .A0(n14374), .A1(n14365), .S(n4165), .Z(n14381) );
  CMX2X1 U25322 ( .A0(n14366), .A1(n14381), .S(n4313), .Z(n14394) );
  CMXI2X1 U25323 ( .A0(n14367), .A1(n14394), .S(n3361), .Z(N8868) );
  CMX2X1 U25324 ( .A0(N7676), .A1(N7675), .S(n3868), .Z(n14377) );
  CMXI2X1 U25325 ( .A0(n14377), .A1(n14368), .S(n4165), .Z(n14384) );
  CMX2X1 U25326 ( .A0(n14369), .A1(n14384), .S(n4312), .Z(n14397) );
  CMXI2X1 U25327 ( .A0(n14370), .A1(n14397), .S(n3361), .Z(N8869) );
  CMX2X1 U25328 ( .A0(N8207), .A1(N8206), .S(n3869), .Z(n14441) );
  CMXI2X1 U25329 ( .A0(n14441), .A1(n14371), .S(n4164), .Z(n14508) );
  CMX2X1 U25330 ( .A0(n14372), .A1(n14508), .S(n4312), .Z(n14641) );
  CMXI2X1 U25331 ( .A0(n14373), .A1(n14641), .S(n3361), .Z(N8338) );
  CMX2X1 U25332 ( .A0(N7675), .A1(N7674), .S(n3870), .Z(n14380) );
  CMXI2X1 U25333 ( .A0(n14380), .A1(n14374), .S(n4164), .Z(n14387) );
  CMX2X1 U25334 ( .A0(n14375), .A1(n14387), .S(n4312), .Z(n14400) );
  CMXI2X1 U25335 ( .A0(n14376), .A1(n14400), .S(n3361), .Z(N8870) );
  CMX2X1 U25336 ( .A0(N7674), .A1(N7673), .S(n3871), .Z(n14383) );
  CMXI2X1 U25337 ( .A0(n14383), .A1(n14377), .S(n4164), .Z(n14390) );
  CMX2X1 U25338 ( .A0(n14378), .A1(n14390), .S(n4312), .Z(n14403) );
  CMXI2X1 U25339 ( .A0(n14379), .A1(n14403), .S(n3361), .Z(N8871) );
  CMX2X1 U25340 ( .A0(N7673), .A1(N7672), .S(n3872), .Z(n14386) );
  CMXI2X1 U25341 ( .A0(n14386), .A1(n14380), .S(n4164), .Z(n14393) );
  CMX2X1 U25342 ( .A0(n14381), .A1(n14393), .S(n4312), .Z(n14413) );
  CMXI2X1 U25343 ( .A0(n14382), .A1(n14413), .S(n3361), .Z(N8872) );
  CMX2X1 U25344 ( .A0(N7672), .A1(N7671), .S(n3873), .Z(n14389) );
  CMXI2X1 U25345 ( .A0(n14389), .A1(n14383), .S(n4164), .Z(n14396) );
  CMX2X1 U25346 ( .A0(n14384), .A1(n14396), .S(n4312), .Z(n14416) );
  CMXI2X1 U25347 ( .A0(n14385), .A1(n14416), .S(n3361), .Z(N8873) );
  CMX2X1 U25348 ( .A0(N7671), .A1(N7670), .S(n3874), .Z(n14392) );
  CMXI2X1 U25349 ( .A0(n14392), .A1(n14386), .S(n4164), .Z(n14399) );
  CMX2X1 U25350 ( .A0(n14387), .A1(n14399), .S(n4312), .Z(n14419) );
  CMXI2X1 U25351 ( .A0(n14388), .A1(n14419), .S(n3360), .Z(N8874) );
  CMX2X1 U25352 ( .A0(N7670), .A1(N7669), .S(n3864), .Z(n14395) );
  CMXI2X1 U25353 ( .A0(n14395), .A1(n14389), .S(n4164), .Z(n14402) );
  CMX2X1 U25354 ( .A0(n14390), .A1(n14402), .S(n4312), .Z(n14422) );
  CMXI2X1 U25355 ( .A0(n14391), .A1(n14422), .S(n3360), .Z(N8875) );
  CMX2X1 U25356 ( .A0(N7669), .A1(N7668), .S(n3865), .Z(n14398) );
  CMXI2X1 U25357 ( .A0(n14398), .A1(n14392), .S(n4164), .Z(n14412) );
  CMX2X1 U25358 ( .A0(n14393), .A1(n14412), .S(n4312), .Z(n14425) );
  CMXI2X1 U25359 ( .A0(n14394), .A1(n14425), .S(n3360), .Z(N8876) );
  CMX2X1 U25360 ( .A0(N7668), .A1(N7667), .S(n3875), .Z(n14401) );
  CMXI2X1 U25361 ( .A0(n14401), .A1(n14395), .S(n4164), .Z(n14415) );
  CMX2X1 U25362 ( .A0(n14396), .A1(n14415), .S(n4312), .Z(n14428) );
  CMXI2X1 U25363 ( .A0(n14397), .A1(n14428), .S(n3360), .Z(N8877) );
  CMX2X1 U25364 ( .A0(N7667), .A1(N7666), .S(n3876), .Z(n14411) );
  CMXI2X1 U25365 ( .A0(n14411), .A1(n14398), .S(n4164), .Z(n14418) );
  CMX2X1 U25366 ( .A0(n14399), .A1(n14418), .S(n4312), .Z(n14431) );
  CMXI2X1 U25367 ( .A0(n14400), .A1(n14431), .S(n3360), .Z(N8878) );
  CMX2X1 U25368 ( .A0(N7666), .A1(N7665), .S(n3873), .Z(n14414) );
  CMXI2X1 U25369 ( .A0(n14414), .A1(n14401), .S(n4164), .Z(n14421) );
  CMX2X1 U25370 ( .A0(n14402), .A1(n14421), .S(n4311), .Z(n14434) );
  CMXI2X1 U25371 ( .A0(n14403), .A1(n14434), .S(n3360), .Z(N8879) );
  CMX2X1 U25372 ( .A0(N8206), .A1(N8205), .S(n3874), .Z(n14474) );
  CMXI2X1 U25373 ( .A0(n14474), .A1(n14404), .S(n4164), .Z(n14541) );
  CMX2X1 U25374 ( .A0(n14405), .A1(n14541), .S(n4311), .Z(n14674) );
  CMXI2X1 U25375 ( .A0(n14406), .A1(n14674), .S(n3360), .Z(N8339) );
  CMXI2X1 U25376 ( .A0(n14410), .A1(n14409), .S(n3360), .Z(N8285) );
  CMX2X1 U25377 ( .A0(N7665), .A1(N7664), .S(n3875), .Z(n14417) );
  CMXI2X1 U25378 ( .A0(n14417), .A1(n14411), .S(n4164), .Z(n14424) );
  CMX2X1 U25379 ( .A0(n14412), .A1(n14424), .S(n4311), .Z(n14437) );
  CMXI2X1 U25380 ( .A0(n14413), .A1(n14437), .S(n3363), .Z(N8880) );
  CMX2X1 U25381 ( .A0(N7664), .A1(N7663), .S(n3876), .Z(n14420) );
  CMXI2X1 U25382 ( .A0(n14420), .A1(n14414), .S(n4164), .Z(n14427) );
  CMX2X1 U25383 ( .A0(n14415), .A1(n14427), .S(n4311), .Z(n14440) );
  CMXI2X1 U25384 ( .A0(n14416), .A1(n14440), .S(n3363), .Z(N8881) );
  CMX2X1 U25385 ( .A0(N7663), .A1(N7662), .S(n3871), .Z(n14423) );
  CMXI2X1 U25386 ( .A0(n14423), .A1(n14417), .S(n4164), .Z(n14430) );
  CMX2X1 U25387 ( .A0(n14418), .A1(n14430), .S(n4311), .Z(n14446) );
  CMXI2X1 U25388 ( .A0(n14419), .A1(n14446), .S(n3363), .Z(N8882) );
  CMX2X1 U25389 ( .A0(N7662), .A1(N7661), .S(n3872), .Z(n14426) );
  CMXI2X1 U25390 ( .A0(n14426), .A1(n14420), .S(n4164), .Z(n14433) );
  CMX2X1 U25391 ( .A0(n14421), .A1(n14433), .S(n4311), .Z(n14449) );
  CMXI2X1 U25392 ( .A0(n14422), .A1(n14449), .S(n3363), .Z(N8883) );
  CMX2X1 U25393 ( .A0(N7661), .A1(N7660), .S(n3873), .Z(n14429) );
  CMXI2X1 U25394 ( .A0(n14429), .A1(n14423), .S(n4163), .Z(n14436) );
  CMX2X1 U25395 ( .A0(n14424), .A1(n14436), .S(n4311), .Z(n14452) );
  CMXI2X1 U25396 ( .A0(n14425), .A1(n14452), .S(n3363), .Z(N8884) );
  CMX2X1 U25397 ( .A0(N7660), .A1(N7659), .S(n3874), .Z(n14432) );
  CMXI2X1 U25398 ( .A0(n14432), .A1(n14426), .S(n4163), .Z(n14439) );
  CMX2X1 U25399 ( .A0(n14427), .A1(n14439), .S(n4311), .Z(n14455) );
  CMXI2X1 U25400 ( .A0(n14428), .A1(n14455), .S(n3363), .Z(N8885) );
  CMX2X1 U25401 ( .A0(N7659), .A1(N7658), .S(n3869), .Z(n14435) );
  CMXI2X1 U25402 ( .A0(n14435), .A1(n14429), .S(n4163), .Z(n14445) );
  CMX2X1 U25403 ( .A0(n14430), .A1(n14445), .S(n4311), .Z(n14458) );
  CMXI2X1 U25404 ( .A0(n14431), .A1(n14458), .S(n3362), .Z(N8886) );
  CMX2X1 U25405 ( .A0(N7658), .A1(N7657), .S(n3877), .Z(n14438) );
  CMXI2X1 U25406 ( .A0(n14438), .A1(n14432), .S(n4163), .Z(n14448) );
  CMX2X1 U25407 ( .A0(n14433), .A1(n14448), .S(n4311), .Z(n14461) );
  CMXI2X1 U25408 ( .A0(n14434), .A1(n14461), .S(n3362), .Z(N8887) );
  CMX2X1 U25409 ( .A0(N7657), .A1(N7656), .S(n3878), .Z(n14444) );
  CMXI2X1 U25410 ( .A0(n14444), .A1(n14435), .S(n4163), .Z(n14451) );
  CMX2X1 U25411 ( .A0(n14436), .A1(n14451), .S(n4311), .Z(n14464) );
  CMXI2X1 U25412 ( .A0(n14437), .A1(n14464), .S(n3362), .Z(N8888) );
  CMX2X1 U25413 ( .A0(N7656), .A1(N7655), .S(n3879), .Z(n14447) );
  CMXI2X1 U25414 ( .A0(n14447), .A1(n14438), .S(n4163), .Z(n14454) );
  CMX2X1 U25415 ( .A0(n14439), .A1(n14454), .S(n4310), .Z(n14467) );
  CMXI2X1 U25416 ( .A0(n14440), .A1(n14467), .S(n3362), .Z(N8889) );
  CMX2X1 U25417 ( .A0(N8205), .A1(N8204), .S(n3880), .Z(n14507) );
  CMXI2X1 U25418 ( .A0(n14507), .A1(n14441), .S(n4163), .Z(n14574) );
  CMX2X1 U25419 ( .A0(n14442), .A1(n14574), .S(n4310), .Z(n14707) );
  CMXI2X1 U25420 ( .A0(n14443), .A1(n14707), .S(n3362), .Z(N8340) );
  CMX2X1 U25421 ( .A0(N7655), .A1(N7654), .S(n3881), .Z(n14450) );
  CMXI2X1 U25422 ( .A0(n14450), .A1(n14444), .S(n4163), .Z(n14457) );
  CMX2X1 U25423 ( .A0(n14445), .A1(n14457), .S(n4310), .Z(n14470) );
  CMXI2X1 U25424 ( .A0(n14446), .A1(n14470), .S(n3362), .Z(N8890) );
  CMX2X1 U25425 ( .A0(N7654), .A1(N7653), .S(n3862), .Z(n14453) );
  CMXI2X1 U25426 ( .A0(n14453), .A1(n14447), .S(n4163), .Z(n14460) );
  CMX2X1 U25427 ( .A0(n14448), .A1(n14460), .S(n4310), .Z(n14473) );
  CMXI2X1 U25428 ( .A0(n14449), .A1(n14473), .S(n3362), .Z(N8891) );
  CMX2X1 U25429 ( .A0(N7653), .A1(N7652), .S(n3863), .Z(n14456) );
  CMXI2X1 U25430 ( .A0(n14456), .A1(n14450), .S(n4163), .Z(n14463) );
  CMX2X1 U25431 ( .A0(n14451), .A1(n14463), .S(n4310), .Z(n14479) );
  CMXI2X1 U25432 ( .A0(n14452), .A1(n14479), .S(n3362), .Z(N8892) );
  CMX2X1 U25433 ( .A0(N7652), .A1(N7651), .S(n3866), .Z(n14459) );
  CMXI2X1 U25434 ( .A0(n14459), .A1(n14453), .S(n4163), .Z(n14466) );
  CMX2X1 U25435 ( .A0(n14454), .A1(n14466), .S(n4310), .Z(n14482) );
  CMXI2X1 U25436 ( .A0(n14455), .A1(n14482), .S(n3362), .Z(N8893) );
  CMX2X1 U25437 ( .A0(N7651), .A1(N7650), .S(n3867), .Z(n14462) );
  CMXI2X1 U25438 ( .A0(n14462), .A1(n14456), .S(n4163), .Z(n14469) );
  CMX2X1 U25439 ( .A0(n14457), .A1(n14469), .S(n4310), .Z(n14485) );
  CMXI2X1 U25440 ( .A0(n14458), .A1(n14485), .S(n3362), .Z(N8894) );
  CMX2X1 U25441 ( .A0(N7650), .A1(N7649), .S(n3864), .Z(n14465) );
  CMXI2X1 U25442 ( .A0(n14465), .A1(n14459), .S(n4163), .Z(n14472) );
  CMX2X1 U25443 ( .A0(n14460), .A1(n14472), .S(n4310), .Z(n14488) );
  CMXI2X1 U25444 ( .A0(n14461), .A1(n14488), .S(n3362), .Z(N8895) );
  CMX2X1 U25445 ( .A0(N7649), .A1(N7648), .S(n3865), .Z(n14468) );
  CMXI2X1 U25446 ( .A0(n14468), .A1(n14462), .S(n4163), .Z(n14478) );
  CMX2X1 U25447 ( .A0(n14463), .A1(n14478), .S(n4310), .Z(n14491) );
  CMXI2X1 U25448 ( .A0(n14464), .A1(n14491), .S(n3361), .Z(N8896) );
  CMX2X1 U25449 ( .A0(N7648), .A1(N7647), .S(n3877), .Z(n14471) );
  CMXI2X1 U25450 ( .A0(n14471), .A1(n14465), .S(n4163), .Z(n14481) );
  CMX2X1 U25451 ( .A0(n14466), .A1(n14481), .S(n4310), .Z(n14494) );
  CMXI2X1 U25452 ( .A0(n14467), .A1(n14494), .S(n3365), .Z(N8897) );
  CMX2X1 U25453 ( .A0(N7647), .A1(N7646), .S(n3878), .Z(n14477) );
  CMXI2X1 U25454 ( .A0(n14477), .A1(n14468), .S(n4163), .Z(n14484) );
  CMX2X1 U25455 ( .A0(n14469), .A1(n14484), .S(n4310), .Z(n14497) );
  CMXI2X1 U25456 ( .A0(n14470), .A1(n14497), .S(n3365), .Z(N8898) );
  CMX2X1 U25457 ( .A0(N7646), .A1(N7645), .S(n3879), .Z(n14480) );
  CMXI2X1 U25458 ( .A0(n14480), .A1(n14471), .S(n4162), .Z(n14487) );
  CMX2X1 U25459 ( .A0(n14472), .A1(n14487), .S(n4309), .Z(n14500) );
  CMXI2X1 U25460 ( .A0(n14473), .A1(n14500), .S(n3364), .Z(N8899) );
  CMX2X1 U25461 ( .A0(N8204), .A1(N8203), .S(n3880), .Z(n14540) );
  CMXI2X1 U25462 ( .A0(n14540), .A1(n14474), .S(n4162), .Z(n14607) );
  CMX2X1 U25463 ( .A0(n14475), .A1(n14607), .S(n4309), .Z(n14740) );
  CMXI2X1 U25464 ( .A0(n14476), .A1(n14740), .S(n3364), .Z(N8341) );
  CMX2X1 U25465 ( .A0(N7645), .A1(N7644), .S(n3875), .Z(n14483) );
  CMXI2X1 U25466 ( .A0(n14483), .A1(n14477), .S(n4162), .Z(n14490) );
  CMX2X1 U25467 ( .A0(n14478), .A1(n14490), .S(n4309), .Z(n14503) );
  CMXI2X1 U25468 ( .A0(n14479), .A1(n14503), .S(n3364), .Z(N8900) );
  CMX2X1 U25469 ( .A0(N7644), .A1(N7643), .S(n3876), .Z(n14486) );
  CMXI2X1 U25470 ( .A0(n14486), .A1(n14480), .S(n4162), .Z(n14493) );
  CMX2X1 U25471 ( .A0(n14481), .A1(n14493), .S(n4309), .Z(n14506) );
  CMXI2X1 U25472 ( .A0(n14482), .A1(n14506), .S(n3364), .Z(N8901) );
  CMX2X1 U25473 ( .A0(N7643), .A1(N7642), .S(n3877), .Z(n14489) );
  CMXI2X1 U25474 ( .A0(n14489), .A1(n14483), .S(n4162), .Z(n14496) );
  CMX2X1 U25475 ( .A0(n14484), .A1(n14496), .S(n4309), .Z(n14512) );
  CMXI2X1 U25476 ( .A0(n14485), .A1(n14512), .S(n3364), .Z(N8902) );
  CMX2X1 U25477 ( .A0(N7642), .A1(N7641), .S(n3878), .Z(n14492) );
  CMXI2X1 U25478 ( .A0(n14492), .A1(n14486), .S(n4162), .Z(n14499) );
  CMX2X1 U25479 ( .A0(n14487), .A1(n14499), .S(n4309), .Z(n14515) );
  CMXI2X1 U25480 ( .A0(n14488), .A1(n14515), .S(n3364), .Z(N8903) );
  CMX2X1 U25481 ( .A0(N7641), .A1(N7640), .S(n3870), .Z(n14495) );
  CMXI2X1 U25482 ( .A0(n14495), .A1(n14489), .S(n4162), .Z(n14502) );
  CMX2X1 U25483 ( .A0(n14490), .A1(n14502), .S(n4309), .Z(n14518) );
  CMXI2X1 U25484 ( .A0(n14491), .A1(n14518), .S(n3364), .Z(N8904) );
  CMX2X1 U25485 ( .A0(N7640), .A1(N7639), .S(n3866), .Z(n14498) );
  CMXI2X1 U25486 ( .A0(n14498), .A1(n14492), .S(n4162), .Z(n14505) );
  CMX2X1 U25487 ( .A0(n14493), .A1(n14505), .S(n4309), .Z(n14521) );
  CMXI2X1 U25488 ( .A0(n14494), .A1(n14521), .S(n3364), .Z(N8905) );
  CMX2X1 U25489 ( .A0(N7639), .A1(N7638), .S(n3867), .Z(n14501) );
  CMXI2X1 U25490 ( .A0(n14501), .A1(n14495), .S(n4162), .Z(n14511) );
  CMX2X1 U25491 ( .A0(n14496), .A1(n14511), .S(n4309), .Z(n14524) );
  CMXI2X1 U25492 ( .A0(n14497), .A1(n14524), .S(n3364), .Z(N8906) );
  CMX2X1 U25493 ( .A0(N7638), .A1(N7637), .S(n3878), .Z(n14504) );
  CMXI2X1 U25494 ( .A0(n14504), .A1(n14498), .S(n4162), .Z(n14514) );
  CMX2X1 U25495 ( .A0(n14499), .A1(n14514), .S(n4309), .Z(n14527) );
  CMXI2X1 U25496 ( .A0(n14500), .A1(n14527), .S(n3364), .Z(N8907) );
  CMX2X1 U25497 ( .A0(N7637), .A1(N7636), .S(n3881), .Z(n14510) );
  CMXI2X1 U25498 ( .A0(n14510), .A1(n14501), .S(n4162), .Z(n14517) );
  CMX2X1 U25499 ( .A0(n14502), .A1(n14517), .S(n4309), .Z(n14530) );
  CMXI2X1 U25500 ( .A0(n14503), .A1(n14530), .S(n3364), .Z(N8908) );
  CMX2X1 U25501 ( .A0(N7636), .A1(N7635), .S(n3862), .Z(n14513) );
  CMXI2X1 U25502 ( .A0(n14513), .A1(n14504), .S(n4162), .Z(n14520) );
  CMX2X1 U25503 ( .A0(n14505), .A1(n14520), .S(n4308), .Z(n14533) );
  CMXI2X1 U25504 ( .A0(n14506), .A1(n14533), .S(n3363), .Z(N8909) );
  CMX2X1 U25505 ( .A0(N8203), .A1(N8202), .S(n3866), .Z(n14573) );
  CMXI2X1 U25506 ( .A0(n14573), .A1(n14507), .S(n4162), .Z(n14640) );
  CMX2X1 U25507 ( .A0(n14508), .A1(n14640), .S(n4308), .Z(n14777) );
  CMXI2X1 U25508 ( .A0(n14509), .A1(n14777), .S(n3363), .Z(N8342) );
  CMX2X1 U25509 ( .A0(N7635), .A1(N7634), .S(n3870), .Z(n14516) );
  CMXI2X1 U25510 ( .A0(n14516), .A1(n14510), .S(n4162), .Z(n14523) );
  CMX2X1 U25511 ( .A0(n14511), .A1(n14523), .S(n4308), .Z(n14536) );
  CMXI2X1 U25512 ( .A0(n14512), .A1(n14536), .S(n3363), .Z(N8910) );
  CMX2X1 U25513 ( .A0(N7634), .A1(N7633), .S(n3871), .Z(n14519) );
  CMXI2X1 U25514 ( .A0(n14519), .A1(n14513), .S(n4162), .Z(n14526) );
  CMX2X1 U25515 ( .A0(n14514), .A1(n14526), .S(n4308), .Z(n14539) );
  CMXI2X1 U25516 ( .A0(n14515), .A1(n14539), .S(n3363), .Z(N8911) );
  CMX2X1 U25517 ( .A0(N7633), .A1(N7632), .S(n3872), .Z(n14522) );
  CMXI2X1 U25518 ( .A0(n14522), .A1(n14516), .S(n4162), .Z(n14529) );
  CMX2X1 U25519 ( .A0(n14517), .A1(n14529), .S(n4308), .Z(n14545) );
  CMXI2X1 U25520 ( .A0(n14518), .A1(n14545), .S(n3363), .Z(N8912) );
  CMX2X1 U25521 ( .A0(N7632), .A1(N7631), .S(n3873), .Z(n14525) );
  CMXI2X1 U25522 ( .A0(n14525), .A1(n14519), .S(n4161), .Z(n14532) );
  CMX2X1 U25523 ( .A0(n14520), .A1(n14532), .S(n4308), .Z(n14548) );
  CMXI2X1 U25524 ( .A0(n14521), .A1(n14548), .S(n3333), .Z(N8913) );
  CMX2X1 U25525 ( .A0(N7631), .A1(N7630), .S(n3874), .Z(n14528) );
  CMXI2X1 U25526 ( .A0(n14528), .A1(n14522), .S(n4161), .Z(n14535) );
  CMX2X1 U25527 ( .A0(n14523), .A1(n14535), .S(n4308), .Z(n14551) );
  CMXI2X1 U25528 ( .A0(n14524), .A1(n14551), .S(n3333), .Z(N8914) );
  CMX2X1 U25529 ( .A0(N7630), .A1(N7629), .S(n3875), .Z(n14531) );
  CMXI2X1 U25530 ( .A0(n14531), .A1(n14525), .S(n4161), .Z(n14538) );
  CMX2X1 U25531 ( .A0(n14526), .A1(n14538), .S(n4308), .Z(n14554) );
  CMXI2X1 U25532 ( .A0(n14527), .A1(n14554), .S(n3333), .Z(N8915) );
  CMX2X1 U25533 ( .A0(N7629), .A1(N7628), .S(n3876), .Z(n14534) );
  CMXI2X1 U25534 ( .A0(n14534), .A1(n14528), .S(n4161), .Z(n14544) );
  CMX2X1 U25535 ( .A0(n14529), .A1(n14544), .S(n4308), .Z(n14557) );
  CMXI2X1 U25536 ( .A0(n14530), .A1(n14557), .S(n3333), .Z(N8916) );
  CMX2X1 U25537 ( .A0(N7628), .A1(N7627), .S(n3880), .Z(n14537) );
  CMXI2X1 U25538 ( .A0(n14537), .A1(n14531), .S(n4161), .Z(n14547) );
  CMX2X1 U25539 ( .A0(n14532), .A1(n14547), .S(n4308), .Z(n14560) );
  CMXI2X1 U25540 ( .A0(n14533), .A1(n14560), .S(n3332), .Z(N8917) );
  CMX2X1 U25541 ( .A0(N7627), .A1(N7626), .S(n3881), .Z(n14543) );
  CMXI2X1 U25542 ( .A0(n14543), .A1(n14534), .S(n4161), .Z(n14550) );
  CMX2X1 U25543 ( .A0(n14535), .A1(n14550), .S(n4308), .Z(n14563) );
  CMXI2X1 U25544 ( .A0(n14536), .A1(n14563), .S(n3332), .Z(N8918) );
  CMX2X1 U25545 ( .A0(N7626), .A1(N7625), .S(n3877), .Z(n14546) );
  CMXI2X1 U25546 ( .A0(n14546), .A1(n14537), .S(n4161), .Z(n14553) );
  CMX2X1 U25547 ( .A0(n14538), .A1(n14553), .S(n4307), .Z(n14566) );
  CMXI2X1 U25548 ( .A0(n14539), .A1(n14566), .S(n3340), .Z(N8919) );
  CMX2X1 U25549 ( .A0(N8202), .A1(N8201), .S(n3878), .Z(n14606) );
  CMXI2X1 U25550 ( .A0(n14606), .A1(n14540), .S(n4161), .Z(n14673) );
  CMX2X1 U25551 ( .A0(n14541), .A1(n14673), .S(n4316), .Z(n14810) );
  CMXI2X1 U25552 ( .A0(n14542), .A1(n14810), .S(n3391), .Z(N8343) );
  CMX2X1 U25553 ( .A0(N7625), .A1(N7624), .S(n3865), .Z(n14549) );
  CMXI2X1 U25554 ( .A0(n14549), .A1(n14543), .S(n4161), .Z(n14556) );
  CMX2X1 U25555 ( .A0(n14544), .A1(n14556), .S(n3776), .Z(n14569) );
  CMXI2X1 U25556 ( .A0(n14545), .A1(n14569), .S(n3356), .Z(N8920) );
  CMX2X1 U25557 ( .A0(N7624), .A1(N7623), .S(n3866), .Z(n14552) );
  CMXI2X1 U25558 ( .A0(n14552), .A1(n14546), .S(n4161), .Z(n14559) );
  CMX2X1 U25559 ( .A0(n14547), .A1(n14559), .S(n3777), .Z(n14572) );
  CMXI2X1 U25560 ( .A0(n14548), .A1(n14572), .S(n3365), .Z(N8921) );
  CMX2X1 U25561 ( .A0(N7623), .A1(N7622), .S(n3867), .Z(n14555) );
  CMXI2X1 U25562 ( .A0(n14555), .A1(n14549), .S(n4161), .Z(n14562) );
  CMX2X1 U25563 ( .A0(n14550), .A1(n14562), .S(n3790), .Z(n14578) );
  CMXI2X1 U25564 ( .A0(n14551), .A1(n14578), .S(n3365), .Z(N8922) );
  CMX2X1 U25565 ( .A0(N7622), .A1(N7621), .S(n3868), .Z(n14558) );
  CMXI2X1 U25566 ( .A0(n14558), .A1(n14552), .S(n4161), .Z(n14565) );
  CMX2X1 U25567 ( .A0(n14553), .A1(n14565), .S(n3791), .Z(n14581) );
  CMXI2X1 U25568 ( .A0(n14554), .A1(n14581), .S(n3365), .Z(N8923) );
  CMX2X1 U25569 ( .A0(N7621), .A1(N7620), .S(n3863), .Z(n14561) );
  CMXI2X1 U25570 ( .A0(n14561), .A1(n14555), .S(n4161), .Z(n14568) );
  CMX2X1 U25571 ( .A0(n14556), .A1(n14568), .S(n3810), .Z(n14584) );
  CMXI2X1 U25572 ( .A0(n14557), .A1(n14584), .S(n3365), .Z(N8924) );
  CMX2X1 U25573 ( .A0(N7620), .A1(N7619), .S(n3864), .Z(n14564) );
  CMXI2X1 U25574 ( .A0(n14564), .A1(n14558), .S(n4161), .Z(n14571) );
  CMX2X1 U25575 ( .A0(n14559), .A1(n14571), .S(n3795), .Z(n14587) );
  CMXI2X1 U25576 ( .A0(n14560), .A1(n14587), .S(n3365), .Z(N8925) );
  CMX2X1 U25577 ( .A0(N7619), .A1(N7618), .S(n3865), .Z(n14567) );
  CMXI2X1 U25578 ( .A0(n14567), .A1(n14561), .S(n4161), .Z(n14577) );
  CMX2X1 U25579 ( .A0(n14562), .A1(n14577), .S(n3811), .Z(n14590) );
  CMXI2X1 U25580 ( .A0(n14563), .A1(n14590), .S(n3365), .Z(N8926) );
  CMX2X1 U25581 ( .A0(N7618), .A1(N7617), .S(n3866), .Z(n14570) );
  CMXI2X1 U25582 ( .A0(n14570), .A1(n14564), .S(n4161), .Z(n14580) );
  CMX2X1 U25583 ( .A0(n14565), .A1(n14580), .S(n3812), .Z(n14593) );
  CMXI2X1 U25584 ( .A0(n14566), .A1(n14593), .S(n3365), .Z(N8927) );
  CMX2X1 U25585 ( .A0(N7617), .A1(N7616), .S(n3867), .Z(n14576) );
  CMXI2X1 U25586 ( .A0(n14576), .A1(n14567), .S(n4160), .Z(n14583) );
  CMX2X1 U25587 ( .A0(n14568), .A1(n14583), .S(n4305), .Z(n14596) );
  CMXI2X1 U25588 ( .A0(n14569), .A1(n14596), .S(n3365), .Z(N8928) );
  CMX2X1 U25589 ( .A0(N7616), .A1(N7615), .S(n3879), .Z(n14579) );
  CMXI2X1 U25590 ( .A0(n14579), .A1(n14570), .S(n4160), .Z(n14586) );
  CMX2X1 U25591 ( .A0(n14571), .A1(n14586), .S(n3771), .Z(n14599) );
  CMXI2X1 U25592 ( .A0(n14572), .A1(n14599), .S(n3365), .Z(N8929) );
  CMX2X1 U25593 ( .A0(N8201), .A1(N8200), .S(n3880), .Z(n14639) );
  CMXI2X1 U25594 ( .A0(n14639), .A1(n14573), .S(n4160), .Z(n14706) );
  CMX2X1 U25595 ( .A0(n14574), .A1(n14706), .S(n3772), .Z(n14843) );
  CMXI2X1 U25596 ( .A0(n14575), .A1(n14843), .S(n3331), .Z(N8344) );
  CMX2X1 U25597 ( .A0(N7615), .A1(N7614), .S(n3881), .Z(n14582) );
  CMXI2X1 U25598 ( .A0(n14582), .A1(n14576), .S(n4160), .Z(n14589) );
  CMX2X1 U25599 ( .A0(n14577), .A1(n14589), .S(n3774), .Z(n14602) );
  CMXI2X1 U25600 ( .A0(n14578), .A1(n14602), .S(n3330), .Z(N8930) );
  CMX2X1 U25601 ( .A0(N7614), .A1(N7613), .S(n3862), .Z(n14585) );
  CMXI2X1 U25602 ( .A0(n14585), .A1(n14579), .S(n4160), .Z(n14592) );
  CMX2X1 U25603 ( .A0(n14580), .A1(n14592), .S(n3792), .Z(n14605) );
  CMXI2X1 U25604 ( .A0(n14581), .A1(n14605), .S(n3329), .Z(N8931) );
  CMX2X1 U25605 ( .A0(N7613), .A1(N7612), .S(n3863), .Z(n14588) );
  CMXI2X1 U25606 ( .A0(n14588), .A1(n14582), .S(n4160), .Z(n14595) );
  CMX2X1 U25607 ( .A0(n14583), .A1(n14595), .S(n3793), .Z(n14611) );
  CMXI2X1 U25608 ( .A0(n14584), .A1(n14611), .S(n3328), .Z(N8932) );
  CMX2X1 U25609 ( .A0(N7612), .A1(N7611), .S(n3864), .Z(n14591) );
  CMXI2X1 U25610 ( .A0(n14591), .A1(n14585), .S(n4160), .Z(n14598) );
  CMX2X1 U25611 ( .A0(n14586), .A1(n14598), .S(n3794), .Z(n14614) );
  CMXI2X1 U25612 ( .A0(n14587), .A1(n14614), .S(n3435), .Z(N8933) );
  CMX2X1 U25613 ( .A0(N7611), .A1(N7610), .S(n3865), .Z(n14594) );
  CMXI2X1 U25614 ( .A0(n14594), .A1(n14588), .S(n4160), .Z(n14601) );
  CMX2X1 U25615 ( .A0(n14589), .A1(n14601), .S(n3795), .Z(n14617) );
  CMXI2X1 U25616 ( .A0(n14590), .A1(n14617), .S(n3434), .Z(N8934) );
  CMX2X1 U25617 ( .A0(N7610), .A1(N7609), .S(n3862), .Z(n14597) );
  CMXI2X1 U25618 ( .A0(n14597), .A1(n14591), .S(n4160), .Z(n14604) );
  CMX2X1 U25619 ( .A0(n14592), .A1(n14604), .S(n3796), .Z(n14620) );
  CMXI2X1 U25620 ( .A0(n14593), .A1(n14620), .S(n3371), .Z(N8935) );
  CMX2X1 U25621 ( .A0(N7609), .A1(N7608), .S(n3863), .Z(n14600) );
  CMXI2X1 U25622 ( .A0(n14600), .A1(n14594), .S(n4160), .Z(n14610) );
  CMX2X1 U25623 ( .A0(n14595), .A1(n14610), .S(n3797), .Z(n14623) );
  CMXI2X1 U25624 ( .A0(n14596), .A1(n14623), .S(n3379), .Z(N8936) );
  CMX2X1 U25625 ( .A0(N7608), .A1(N7607), .S(n3866), .Z(n14603) );
  CMXI2X1 U25626 ( .A0(n14603), .A1(n14597), .S(n4160), .Z(n14613) );
  CMX2X1 U25627 ( .A0(n14598), .A1(n14613), .S(n3805), .Z(n14626) );
  CMXI2X1 U25628 ( .A0(n14599), .A1(n14626), .S(n3372), .Z(N8937) );
  CMX2X1 U25629 ( .A0(N7607), .A1(N7606), .S(n3867), .Z(n14609) );
  CMXI2X1 U25630 ( .A0(n14609), .A1(n14600), .S(n4160), .Z(n14616) );
  CMX2X1 U25631 ( .A0(n14601), .A1(n14616), .S(n3806), .Z(n14629) );
  CMXI2X1 U25632 ( .A0(n14602), .A1(n14629), .S(n3394), .Z(N8938) );
  CMX2X1 U25633 ( .A0(N7606), .A1(N7605), .S(n3869), .Z(n14612) );
  CMXI2X1 U25634 ( .A0(n14612), .A1(n14603), .S(n4160), .Z(n14619) );
  CMX2X1 U25635 ( .A0(n14604), .A1(n14619), .S(n3807), .Z(n14632) );
  CMXI2X1 U25636 ( .A0(n14605), .A1(n14632), .S(n3394), .Z(N8939) );
  CMX2X1 U25637 ( .A0(N8200), .A1(N8199), .S(n3870), .Z(n14672) );
  CMXI2X1 U25638 ( .A0(n14672), .A1(n14606), .S(n4160), .Z(n14739) );
  CMX2X1 U25639 ( .A0(n14607), .A1(n14739), .S(n3808), .Z(n14876) );
  CMXI2X1 U25640 ( .A0(n14608), .A1(n14876), .S(n3394), .Z(N8345) );
  CMX2X1 U25641 ( .A0(N7605), .A1(N7604), .S(n3871), .Z(n14615) );
  CMXI2X1 U25642 ( .A0(n14615), .A1(n14609), .S(n4160), .Z(n14622) );
  CMX2X1 U25643 ( .A0(n14610), .A1(n14622), .S(n3809), .Z(n14635) );
  CMXI2X1 U25644 ( .A0(n14611), .A1(n14635), .S(n3394), .Z(N8940) );
  CMX2X1 U25645 ( .A0(N7604), .A1(N7603), .S(n3872), .Z(n14618) );
  CMXI2X1 U25646 ( .A0(n14618), .A1(n14612), .S(n4160), .Z(n14625) );
  CMX2X1 U25647 ( .A0(n14613), .A1(n14625), .S(n3810), .Z(n14638) );
  CMXI2X1 U25648 ( .A0(n14614), .A1(n14638), .S(n3394), .Z(N8941) );
  CMX2X1 U25649 ( .A0(N7603), .A1(N7602), .S(n3867), .Z(n14621) );
  CMXI2X1 U25650 ( .A0(n14621), .A1(n14615), .S(n4159), .Z(n14628) );
  CMX2X1 U25651 ( .A0(n14616), .A1(n14628), .S(n3811), .Z(n14644) );
  CMXI2X1 U25652 ( .A0(n14617), .A1(n14644), .S(n3366), .Z(N8942) );
  CMX2X1 U25653 ( .A0(N7602), .A1(N7601), .S(n3868), .Z(n14624) );
  CMXI2X1 U25654 ( .A0(n14624), .A1(n14618), .S(n4159), .Z(n14631) );
  CMX2X1 U25655 ( .A0(n14619), .A1(n14631), .S(n3812), .Z(n14647) );
  CMXI2X1 U25656 ( .A0(n14620), .A1(n14647), .S(n3366), .Z(N8943) );
  CMX2X1 U25657 ( .A0(N7601), .A1(N7600), .S(n3869), .Z(n14627) );
  CMXI2X1 U25658 ( .A0(n14627), .A1(n14621), .S(n4159), .Z(n14634) );
  CMX2X1 U25659 ( .A0(n14622), .A1(n14634), .S(n4305), .Z(n14650) );
  CMXI2X1 U25660 ( .A0(n14623), .A1(n14650), .S(n3366), .Z(N8944) );
  CMX2X1 U25661 ( .A0(N7600), .A1(N7599), .S(n3870), .Z(n14630) );
  CMXI2X1 U25662 ( .A0(n14630), .A1(n14624), .S(n4159), .Z(n14637) );
  CMX2X1 U25663 ( .A0(n14625), .A1(n14637), .S(n3771), .Z(n14653) );
  CMXI2X1 U25664 ( .A0(n14626), .A1(n14653), .S(n3366), .Z(N8945) );
  CMX2X1 U25665 ( .A0(N7599), .A1(N7598), .S(n3868), .Z(n14633) );
  CMXI2X1 U25666 ( .A0(n14633), .A1(n14627), .S(n4159), .Z(n14643) );
  CMX2X1 U25667 ( .A0(n14628), .A1(n14643), .S(n3811), .Z(n14656) );
  CMXI2X1 U25668 ( .A0(n14629), .A1(n14656), .S(n3366), .Z(N8946) );
  CMX2X1 U25669 ( .A0(N7598), .A1(N7597), .S(n3868), .Z(n14636) );
  CMXI2X1 U25670 ( .A0(n14636), .A1(n14630), .S(n4159), .Z(n14646) );
  CMX2X1 U25671 ( .A0(n14631), .A1(n14646), .S(n3796), .Z(n14659) );
  CMXI2X1 U25672 ( .A0(n14632), .A1(n14659), .S(n3366), .Z(N8947) );
  CMX2X1 U25673 ( .A0(N7597), .A1(N7596), .S(n3869), .Z(n14642) );
  CMXI2X1 U25674 ( .A0(n14642), .A1(n14633), .S(n4159), .Z(n14649) );
  CMX2X1 U25675 ( .A0(n14634), .A1(n14649), .S(n3773), .Z(n14662) );
  CMXI2X1 U25676 ( .A0(n14635), .A1(n14662), .S(n3366), .Z(N8948) );
  CMX2X1 U25677 ( .A0(N7596), .A1(N7595), .S(n3870), .Z(n14645) );
  CMXI2X1 U25678 ( .A0(n14645), .A1(n14636), .S(n4159), .Z(n14652) );
  CMX2X1 U25679 ( .A0(n14637), .A1(n14652), .S(n3774), .Z(n14665) );
  CMXI2X1 U25680 ( .A0(n14638), .A1(n14665), .S(n3366), .Z(N8949) );
  CMX2X1 U25681 ( .A0(N8199), .A1(N8198), .S(n3871), .Z(n14705) );
  CMXI2X1 U25682 ( .A0(n14705), .A1(n14639), .S(n4159), .Z(n14776) );
  CMX2X1 U25683 ( .A0(n14640), .A1(n14776), .S(n3775), .Z(n14909) );
  CMXI2X1 U25684 ( .A0(n14641), .A1(n14909), .S(n3366), .Z(N8346) );
  CMX2X1 U25685 ( .A0(N7595), .A1(N7594), .S(n3872), .Z(n14648) );
  CMXI2X1 U25686 ( .A0(n14648), .A1(n14642), .S(n4159), .Z(n14655) );
  CMX2X1 U25687 ( .A0(n14643), .A1(n14655), .S(n3776), .Z(n14668) );
  CMXI2X1 U25688 ( .A0(n14644), .A1(n14668), .S(n3366), .Z(N8950) );
  CMX2X1 U25689 ( .A0(N7594), .A1(N7593), .S(n3873), .Z(n14651) );
  CMXI2X1 U25690 ( .A0(n14651), .A1(n14645), .S(n4159), .Z(n14658) );
  CMX2X1 U25691 ( .A0(n14646), .A1(n14658), .S(n3777), .Z(n14671) );
  CMXI2X1 U25692 ( .A0(n14647), .A1(n14671), .S(n3366), .Z(N8951) );
  CMX2X1 U25693 ( .A0(N7593), .A1(N7592), .S(n3874), .Z(n14654) );
  CMXI2X1 U25694 ( .A0(n14654), .A1(n14648), .S(n4159), .Z(n14661) );
  CMX2X1 U25695 ( .A0(n14649), .A1(n14661), .S(n3775), .Z(n14677) );
  CMXI2X1 U25696 ( .A0(n14650), .A1(n14677), .S(n3388), .Z(N8952) );
  CMX2X1 U25697 ( .A0(N7592), .A1(N7591), .S(n3864), .Z(n14657) );
  CMXI2X1 U25698 ( .A0(n14657), .A1(n14651), .S(n4159), .Z(n14664) );
  CMX2X1 U25699 ( .A0(n14652), .A1(n14664), .S(n3772), .Z(n14680) );
  CMXI2X1 U25700 ( .A0(n14653), .A1(n14680), .S(n3387), .Z(N8953) );
  CMX2X1 U25701 ( .A0(N7591), .A1(N7590), .S(n3865), .Z(n14660) );
  CMXI2X1 U25702 ( .A0(n14660), .A1(n14654), .S(n4159), .Z(n14667) );
  CMX2X1 U25703 ( .A0(n14655), .A1(n14667), .S(n3773), .Z(n14683) );
  CMXI2X1 U25704 ( .A0(n14656), .A1(n14683), .S(n3386), .Z(N8954) );
  CMX2X1 U25705 ( .A0(N7590), .A1(N7589), .S(n3875), .Z(n14663) );
  CMXI2X1 U25706 ( .A0(n14663), .A1(n14657), .S(n4159), .Z(n14670) );
  CMX2X1 U25707 ( .A0(n14658), .A1(n14670), .S(n3774), .Z(n14686) );
  CMXI2X1 U25708 ( .A0(n14659), .A1(n14686), .S(n3385), .Z(N8955) );
  CMX2X1 U25709 ( .A0(N7589), .A1(N7588), .S(n3873), .Z(n14666) );
  CMXI2X1 U25710 ( .A0(n14666), .A1(n14660), .S(n4159), .Z(n14676) );
  CMX2X1 U25711 ( .A0(n14661), .A1(n14676), .S(n3775), .Z(n14689) );
  CMXI2X1 U25712 ( .A0(n14662), .A1(n14689), .S(n3384), .Z(N8956) );
  CMX2X1 U25713 ( .A0(N7588), .A1(N7587), .S(n3874), .Z(n14669) );
  CMXI2X1 U25714 ( .A0(n14669), .A1(n14663), .S(n4158), .Z(n14679) );
  CMX2X1 U25715 ( .A0(n14664), .A1(n14679), .S(n3776), .Z(n14692) );
  CMXI2X1 U25716 ( .A0(n14665), .A1(n14692), .S(n3383), .Z(N8957) );
  CMX2X1 U25717 ( .A0(N7587), .A1(N7586), .S(n3875), .Z(n14675) );
  CMXI2X1 U25718 ( .A0(n14675), .A1(n14666), .S(n4158), .Z(n14682) );
  CMX2X1 U25719 ( .A0(n14667), .A1(n14682), .S(n3777), .Z(n14695) );
  CMXI2X1 U25720 ( .A0(n14668), .A1(n14695), .S(n3381), .Z(N8958) );
  CMX2X1 U25721 ( .A0(N7586), .A1(N7585), .S(n3876), .Z(n14678) );
  CMXI2X1 U25722 ( .A0(n14678), .A1(n14669), .S(n4158), .Z(n14685) );
  CMX2X1 U25723 ( .A0(n14670), .A1(n14685), .S(n3790), .Z(n14698) );
  CMXI2X1 U25724 ( .A0(n14671), .A1(n14698), .S(n3368), .Z(N8959) );
  CMX2X1 U25725 ( .A0(N8198), .A1(N8197), .S(n3877), .Z(n14738) );
  CMXI2X1 U25726 ( .A0(n14738), .A1(n14672), .S(n4158), .Z(n14809) );
  CMX2X1 U25727 ( .A0(n14673), .A1(n14809), .S(n3791), .Z(n14942) );
  CMXI2X1 U25728 ( .A0(n14674), .A1(n14942), .S(n3368), .Z(N8347) );
  CMX2X1 U25729 ( .A0(N7585), .A1(N7584), .S(n3878), .Z(n14681) );
  CMXI2X1 U25730 ( .A0(n14681), .A1(n14675), .S(n4158), .Z(n14688) );
  CMX2X1 U25731 ( .A0(n14676), .A1(n14688), .S(n3792), .Z(n14701) );
  CMXI2X1 U25732 ( .A0(n14677), .A1(n14701), .S(n3368), .Z(N8960) );
  CMX2X1 U25733 ( .A0(N7584), .A1(N7583), .S(n3879), .Z(n14684) );
  CMXI2X1 U25734 ( .A0(n14684), .A1(n14678), .S(n4158), .Z(n14691) );
  CMX2X1 U25735 ( .A0(n14679), .A1(n14691), .S(n3793), .Z(n14704) );
  CMXI2X1 U25736 ( .A0(n14680), .A1(n14704), .S(n3368), .Z(N8961) );
  CMX2X1 U25737 ( .A0(N7583), .A1(N7582), .S(n3873), .Z(n14687) );
  CMXI2X1 U25738 ( .A0(n14687), .A1(n14681), .S(n4158), .Z(n14694) );
  CMX2X1 U25739 ( .A0(n14682), .A1(n14694), .S(n3794), .Z(n14710) );
  CMXI2X1 U25740 ( .A0(n14683), .A1(n14710), .S(n3368), .Z(N8962) );
  CMX2X1 U25741 ( .A0(N7582), .A1(N7581), .S(n3874), .Z(n14690) );
  CMXI2X1 U25742 ( .A0(n14690), .A1(n14684), .S(n4158), .Z(n14697) );
  CMX2X1 U25743 ( .A0(n14685), .A1(n14697), .S(n3795), .Z(n14713) );
  CMXI2X1 U25744 ( .A0(n14686), .A1(n14713), .S(n3368), .Z(N8963) );
  CMX2X1 U25745 ( .A0(N7581), .A1(N7580), .S(n3880), .Z(n14693) );
  CMXI2X1 U25746 ( .A0(n14693), .A1(n14687), .S(n4158), .Z(n14700) );
  CMX2X1 U25747 ( .A0(n14688), .A1(n14700), .S(n3796), .Z(n14716) );
  CMXI2X1 U25748 ( .A0(n14689), .A1(n14716), .S(n3368), .Z(N8964) );
  CMX2X1 U25749 ( .A0(N7580), .A1(N7579), .S(n3881), .Z(n14696) );
  CMXI2X1 U25750 ( .A0(n14696), .A1(n14690), .S(n4158), .Z(n14703) );
  CMX2X1 U25751 ( .A0(n14691), .A1(n14703), .S(n3797), .Z(n14719) );
  CMXI2X1 U25752 ( .A0(n14692), .A1(n14719), .S(n3367), .Z(N8965) );
  CMX2X1 U25753 ( .A0(N7579), .A1(N7578), .S(n3877), .Z(n14699) );
  CMXI2X1 U25754 ( .A0(n14699), .A1(n14693), .S(n4158), .Z(n14709) );
  CMX2X1 U25755 ( .A0(n14694), .A1(n14709), .S(n3805), .Z(n14722) );
  CMXI2X1 U25756 ( .A0(n14695), .A1(n14722), .S(n3367), .Z(N8966) );
  CMX2X1 U25757 ( .A0(N7578), .A1(N7577), .S(n3878), .Z(n14702) );
  CMXI2X1 U25758 ( .A0(n14702), .A1(n14696), .S(n4158), .Z(n14712) );
  CMX2X1 U25759 ( .A0(n14697), .A1(n14712), .S(n3806), .Z(n14725) );
  CMXI2X1 U25760 ( .A0(n14698), .A1(n14725), .S(n3367), .Z(N8967) );
  CMX2X1 U25761 ( .A0(N7577), .A1(N7576), .S(n3879), .Z(n14708) );
  CMXI2X1 U25762 ( .A0(n14708), .A1(n14699), .S(n4158), .Z(n14715) );
  CMX2X1 U25763 ( .A0(n14700), .A1(n14715), .S(n3812), .Z(n14728) );
  CMXI2X1 U25764 ( .A0(n14701), .A1(n14728), .S(n3367), .Z(N8968) );
  CMX2X1 U25765 ( .A0(N7576), .A1(N7575), .S(n3880), .Z(n14711) );
  CMXI2X1 U25766 ( .A0(n14711), .A1(n14702), .S(n4158), .Z(n14718) );
  CMX2X1 U25767 ( .A0(n14703), .A1(n14718), .S(n3797), .Z(n14731) );
  CMXI2X1 U25768 ( .A0(n14704), .A1(n14731), .S(n3367), .Z(N8969) );
  CMX2X1 U25769 ( .A0(N8197), .A1(N8196), .S(n3870), .Z(n14775) );
  CMXI2X1 U25770 ( .A0(n14775), .A1(n14705), .S(n4158), .Z(n14842) );
  CMX2X1 U25771 ( .A0(n14706), .A1(n14842), .S(n3790), .Z(n14975) );
  CMXI2X1 U25772 ( .A0(n14707), .A1(n14975), .S(n3367), .Z(N8348) );
  CMX2X1 U25773 ( .A0(N7575), .A1(N7574), .S(n3871), .Z(n14714) );
  CMXI2X1 U25774 ( .A0(n14714), .A1(n14708), .S(n4158), .Z(n14721) );
  CMX2X1 U25775 ( .A0(n14709), .A1(n14721), .S(n3791), .Z(n14734) );
  CMXI2X1 U25776 ( .A0(n14710), .A1(n14734), .S(n3367), .Z(N8970) );
  CMX2X1 U25777 ( .A0(N7574), .A1(N7573), .S(n3872), .Z(n14717) );
  CMXI2X1 U25778 ( .A0(n14717), .A1(n14711), .S(n4157), .Z(n14724) );
  CMX2X1 U25779 ( .A0(n14712), .A1(n14724), .S(n3792), .Z(n14737) );
  CMXI2X1 U25780 ( .A0(n14713), .A1(n14737), .S(n3367), .Z(N8971) );
  CMX2X1 U25781 ( .A0(N7573), .A1(N7572), .S(n3873), .Z(n14720) );
  CMXI2X1 U25782 ( .A0(n14720), .A1(n14714), .S(n4157), .Z(n14727) );
  CMX2X1 U25783 ( .A0(n14715), .A1(n14727), .S(n3793), .Z(n14747) );
  CMXI2X1 U25784 ( .A0(n14716), .A1(n14747), .S(n3367), .Z(N8972) );
  CMX2X1 U25785 ( .A0(N7572), .A1(N7571), .S(n3868), .Z(n14723) );
  CMXI2X1 U25786 ( .A0(n14723), .A1(n14717), .S(n4157), .Z(n14730) );
  CMX2X1 U25787 ( .A0(n14718), .A1(n14730), .S(n3794), .Z(n14750) );
  CMXI2X1 U25788 ( .A0(n14719), .A1(n14750), .S(n3367), .Z(N8973) );
  CMX2X1 U25789 ( .A0(N7571), .A1(N7570), .S(n3862), .Z(n14726) );
  CMXI2X1 U25790 ( .A0(n14726), .A1(n14720), .S(n4157), .Z(n14733) );
  CMX2X1 U25791 ( .A0(n14721), .A1(n14733), .S(n3776), .Z(n14753) );
  CMXI2X1 U25792 ( .A0(n14722), .A1(n14753), .S(n3367), .Z(N8974) );
  CMX2X1 U25793 ( .A0(N7570), .A1(N7569), .S(n3863), .Z(n14729) );
  CMXI2X1 U25794 ( .A0(n14729), .A1(n14723), .S(n4157), .Z(n14736) );
  CMX2X1 U25795 ( .A0(n14724), .A1(n14736), .S(n3807), .Z(n14756) );
  CMXI2X1 U25796 ( .A0(n14725), .A1(n14756), .S(n3370), .Z(N8975) );
  CMX2X1 U25797 ( .A0(N7569), .A1(N7568), .S(n3876), .Z(n14732) );
  CMXI2X1 U25798 ( .A0(n14732), .A1(n14726), .S(n4157), .Z(n14746) );
  CMX2X1 U25799 ( .A0(n14727), .A1(n14746), .S(n3808), .Z(n14759) );
  CMXI2X1 U25800 ( .A0(n14728), .A1(n14759), .S(n3370), .Z(N8976) );
  CMX2X1 U25801 ( .A0(N7568), .A1(N7567), .S(n3873), .Z(n14735) );
  CMXI2X1 U25802 ( .A0(n14735), .A1(n14729), .S(n4157), .Z(n14749) );
  CMX2X1 U25803 ( .A0(n14730), .A1(n14749), .S(n3809), .Z(n14762) );
  CMXI2X1 U25804 ( .A0(n14731), .A1(n14762), .S(n3370), .Z(N8977) );
  CMX2X1 U25805 ( .A0(N7567), .A1(N7566), .S(n3874), .Z(n14745) );
  CMXI2X1 U25806 ( .A0(n14745), .A1(n14732), .S(n4157), .Z(n14752) );
  CMX2X1 U25807 ( .A0(n14733), .A1(n14752), .S(n3810), .Z(n14765) );
  CMXI2X1 U25808 ( .A0(n14734), .A1(n14765), .S(n3369), .Z(N8978) );
  CMX2X1 U25809 ( .A0(N7566), .A1(N7565), .S(n3875), .Z(n14748) );
  CMXI2X1 U25810 ( .A0(n14748), .A1(n14735), .S(n4157), .Z(n14755) );
  CMX2X1 U25811 ( .A0(n14736), .A1(n14755), .S(n3811), .Z(n14768) );
  CMXI2X1 U25812 ( .A0(n14737), .A1(n14768), .S(n3369), .Z(N8979) );
  CMX2X1 U25813 ( .A0(N8196), .A1(N8195), .S(n3876), .Z(n14808) );
  CMXI2X1 U25814 ( .A0(n14808), .A1(n14738), .S(n4157), .Z(n14875) );
  CMX2X1 U25815 ( .A0(n14739), .A1(n14875), .S(n3812), .Z(n15008) );
  CMXI2X1 U25816 ( .A0(n14740), .A1(n15008), .S(n3369), .Z(N8349) );
  CMXI2X1 U25817 ( .A0(n4425), .A1(n14742), .S(n3779), .Z(n14744) );
  CMXI2X1 U25818 ( .A0(n14744), .A1(n14743), .S(n3369), .Z(N8286) );
  CMX2X1 U25819 ( .A0(N7565), .A1(N7564), .S(n3871), .Z(n14751) );
  CMXI2X1 U25820 ( .A0(n14751), .A1(n14745), .S(n4157), .Z(n14758) );
  CMX2X1 U25821 ( .A0(n14746), .A1(n14758), .S(n4306), .Z(n14771) );
  CMXI2X1 U25822 ( .A0(n14747), .A1(n14771), .S(n3369), .Z(N8980) );
  CMX2X1 U25823 ( .A0(N7564), .A1(N7563), .S(n3872), .Z(n14754) );
  CMXI2X1 U25824 ( .A0(n14754), .A1(n14748), .S(n4157), .Z(n14761) );
  CMX2X1 U25825 ( .A0(n14749), .A1(n14761), .S(n3771), .Z(n14774) );
  CMXI2X1 U25826 ( .A0(n14750), .A1(n14774), .S(n3369), .Z(N8981) );
  CMX2X1 U25827 ( .A0(N7563), .A1(N7562), .S(n3873), .Z(n14757) );
  CMXI2X1 U25828 ( .A0(n14757), .A1(n14751), .S(n4157), .Z(n14764) );
  CMX2X1 U25829 ( .A0(n14752), .A1(n14764), .S(n3772), .Z(n14780) );
  CMXI2X1 U25830 ( .A0(n14753), .A1(n14780), .S(n3369), .Z(N8982) );
  CMX2X1 U25831 ( .A0(N7562), .A1(N7561), .S(n3874), .Z(n14760) );
  CMXI2X1 U25832 ( .A0(n14760), .A1(n14754), .S(n4157), .Z(n14767) );
  CMX2X1 U25833 ( .A0(n14755), .A1(n14767), .S(n3773), .Z(n14783) );
  CMXI2X1 U25834 ( .A0(n14756), .A1(n14783), .S(n3369), .Z(N8983) );
  CMX2X1 U25835 ( .A0(N7561), .A1(N7560), .S(n3869), .Z(n14763) );
  CMXI2X1 U25836 ( .A0(n14763), .A1(n14757), .S(n4157), .Z(n14770) );
  CMX2X1 U25837 ( .A0(n14758), .A1(n14770), .S(n3774), .Z(n14786) );
  CMXI2X1 U25838 ( .A0(n14759), .A1(n14786), .S(n3369), .Z(N8984) );
  CMX2X1 U25839 ( .A0(N7560), .A1(N7559), .S(n3877), .Z(n14766) );
  CMXI2X1 U25840 ( .A0(n14766), .A1(n14760), .S(n4157), .Z(n14773) );
  CMX2X1 U25841 ( .A0(n14761), .A1(n14773), .S(n3775), .Z(n14789) );
  CMXI2X1 U25842 ( .A0(n14762), .A1(n14789), .S(n3369), .Z(N8985) );
  CMX2X1 U25843 ( .A0(N7559), .A1(N7558), .S(n3878), .Z(n14769) );
  CMXI2X1 U25844 ( .A0(n14769), .A1(n14763), .S(n4156), .Z(n14779) );
  CMX2X1 U25845 ( .A0(n14764), .A1(n14779), .S(n3776), .Z(n14792) );
  CMXI2X1 U25846 ( .A0(n14765), .A1(n14792), .S(n3369), .Z(N8986) );
  CMX2X1 U25847 ( .A0(N7558), .A1(N7557), .S(n3879), .Z(n14772) );
  CMXI2X1 U25848 ( .A0(n14772), .A1(n14766), .S(n4156), .Z(n14782) );
  CMX2X1 U25849 ( .A0(n14767), .A1(n14782), .S(n3777), .Z(n14795) );
  CMXI2X1 U25850 ( .A0(n14768), .A1(n14795), .S(n3368), .Z(N8987) );
  CMX2X1 U25851 ( .A0(N7557), .A1(N7556), .S(n3880), .Z(n14778) );
  CMXI2X1 U25852 ( .A0(n14778), .A1(n14769), .S(n4156), .Z(n14785) );
  CMX2X1 U25853 ( .A0(n14770), .A1(n14785), .S(n3790), .Z(n14798) );
  CMXI2X1 U25854 ( .A0(n14771), .A1(n14798), .S(n3368), .Z(N8988) );
  CMX2X1 U25855 ( .A0(N7556), .A1(N7555), .S(n3881), .Z(n14781) );
  CMXI2X1 U25856 ( .A0(n14781), .A1(n14772), .S(n4156), .Z(n14788) );
  CMX2X1 U25857 ( .A0(n14773), .A1(n14788), .S(n3791), .Z(n14801) );
  CMXI2X1 U25858 ( .A0(n14774), .A1(n14801), .S(n3368), .Z(N8989) );
  CMX2X1 U25859 ( .A0(N8195), .A1(N8194), .S(n3862), .Z(n14841) );
  CMXI2X1 U25860 ( .A0(n14841), .A1(n14775), .S(n4156), .Z(n14908) );
  CMX2X1 U25861 ( .A0(n14776), .A1(n14908), .S(n4306), .Z(n15041) );
  CMXI2X1 U25862 ( .A0(n14777), .A1(n15041), .S(n3368), .Z(N8350) );
  CMX2X1 U25863 ( .A0(N7555), .A1(N7554), .S(n3863), .Z(n14784) );
  CMXI2X1 U25864 ( .A0(n14784), .A1(n14778), .S(n4156), .Z(n14791) );
  CMX2X1 U25865 ( .A0(n14779), .A1(n14791), .S(n3805), .Z(n14804) );
  CMXI2X1 U25866 ( .A0(n14780), .A1(n14804), .S(n3371), .Z(N8990) );
  CMX2X1 U25867 ( .A0(N7554), .A1(N7553), .S(n3866), .Z(n14787) );
  CMXI2X1 U25868 ( .A0(n14787), .A1(n14781), .S(n4156), .Z(n14794) );
  CMX2X1 U25869 ( .A0(n14782), .A1(n14794), .S(n3795), .Z(n14807) );
  CMXI2X1 U25870 ( .A0(n14783), .A1(n14807), .S(n3371), .Z(N8991) );
  CMX2X1 U25871 ( .A0(N7553), .A1(N7552), .S(n3867), .Z(n14790) );
  CMXI2X1 U25872 ( .A0(n14790), .A1(n14784), .S(n4156), .Z(n14797) );
  CMX2X1 U25873 ( .A0(n14785), .A1(n14797), .S(n3796), .Z(n14813) );
  CMXI2X1 U25874 ( .A0(n14786), .A1(n14813), .S(n3371), .Z(N8992) );
  CMX2X1 U25875 ( .A0(N7552), .A1(N7551), .S(n3864), .Z(n14793) );
  CMXI2X1 U25876 ( .A0(n14793), .A1(n14787), .S(n4156), .Z(n14800) );
  CMX2X1 U25877 ( .A0(n14788), .A1(n14800), .S(n3797), .Z(n14816) );
  CMXI2X1 U25878 ( .A0(n14789), .A1(n14816), .S(n3371), .Z(N8993) );
  CMX2X1 U25879 ( .A0(N7551), .A1(N7550), .S(n3877), .Z(n14796) );
  CMXI2X1 U25880 ( .A0(n14796), .A1(n14790), .S(n4156), .Z(n14803) );
  CMX2X1 U25881 ( .A0(n14791), .A1(n14803), .S(n3805), .Z(n14819) );
  CMXI2X1 U25882 ( .A0(n14792), .A1(n14819), .S(n3371), .Z(N8994) );
  CMX2X1 U25883 ( .A0(N7550), .A1(N7549), .S(n3878), .Z(n14799) );
  CMXI2X1 U25884 ( .A0(n14799), .A1(n14793), .S(n4156), .Z(n14806) );
  CMX2X1 U25885 ( .A0(n14794), .A1(n14806), .S(n3806), .Z(n14822) );
  CMXI2X1 U25886 ( .A0(n14795), .A1(n14822), .S(n3371), .Z(N8995) );
  CMX2X1 U25887 ( .A0(N7549), .A1(N7548), .S(n3879), .Z(n14802) );
  CMXI2X1 U25888 ( .A0(n14802), .A1(n14796), .S(n4156), .Z(n14812) );
  CMX2X1 U25889 ( .A0(n14797), .A1(n14812), .S(n3777), .Z(n14825) );
  CMXI2X1 U25890 ( .A0(n14798), .A1(n14825), .S(n3371), .Z(N8996) );
  CMX2X1 U25891 ( .A0(N7548), .A1(N7547), .S(n3880), .Z(n14805) );
  CMXI2X1 U25892 ( .A0(n14805), .A1(n14799), .S(n4156), .Z(n14815) );
  CMX2X1 U25893 ( .A0(n14800), .A1(n14815), .S(n3792), .Z(n14828) );
  CMXI2X1 U25894 ( .A0(n14801), .A1(n14828), .S(n3371), .Z(N8997) );
  CMX2X1 U25895 ( .A0(N7547), .A1(N7546), .S(n3875), .Z(n14811) );
  CMXI2X1 U25896 ( .A0(n14811), .A1(n14802), .S(n4156), .Z(n14818) );
  CMX2X1 U25897 ( .A0(n14803), .A1(n14818), .S(n3793), .Z(n14831) );
  CMXI2X1 U25898 ( .A0(n14804), .A1(n14831), .S(n3371), .Z(N8998) );
  CMX2X1 U25899 ( .A0(N7546), .A1(N7545), .S(n3876), .Z(n14814) );
  CMXI2X1 U25900 ( .A0(n14814), .A1(n14805), .S(n4156), .Z(n14821) );
  CMX2X1 U25901 ( .A0(n14806), .A1(n14821), .S(n3794), .Z(n14834) );
  CMXI2X1 U25902 ( .A0(n14807), .A1(n14834), .S(n3371), .Z(N8999) );
  CMX2X1 U25903 ( .A0(N8194), .A1(N8193), .S(n3877), .Z(n14874) );
  CMXI2X1 U25904 ( .A0(n14874), .A1(n14808), .S(n4156), .Z(n14941) );
  CMX2X1 U25905 ( .A0(n14809), .A1(n14941), .S(n3795), .Z(n15074) );
  CMXI2X1 U25906 ( .A0(n14810), .A1(n15074), .S(n3370), .Z(N8351) );
  CMX2X1 U25907 ( .A0(N7545), .A1(N7544), .S(n3878), .Z(n14817) );
  CMXI2X1 U25908 ( .A0(n14817), .A1(n14811), .S(n4155), .Z(n14824) );
  CMX2X1 U25909 ( .A0(n14812), .A1(n14824), .S(n3796), .Z(n14837) );
  CMXI2X1 U25910 ( .A0(n14813), .A1(n14837), .S(n3370), .Z(N9000) );
  CMX2X1 U25911 ( .A0(N7544), .A1(N7543), .S(n3870), .Z(n14820) );
  CMXI2X1 U25912 ( .A0(n14820), .A1(n14814), .S(n4155), .Z(n14827) );
  CMX2X1 U25913 ( .A0(n14815), .A1(n14827), .S(n3797), .Z(n14840) );
  CMXI2X1 U25914 ( .A0(n14816), .A1(n14840), .S(n3370), .Z(N9001) );
  CMX2X1 U25915 ( .A0(N7543), .A1(N7542), .S(n3866), .Z(n14823) );
  CMXI2X1 U25916 ( .A0(n14823), .A1(n14817), .S(n4155), .Z(n14830) );
  CMX2X1 U25917 ( .A0(n14818), .A1(n14830), .S(n3805), .Z(n14846) );
  CMXI2X1 U25918 ( .A0(n14819), .A1(n14846), .S(n3370), .Z(N9002) );
  CMX2X1 U25919 ( .A0(N7542), .A1(N7541), .S(n3867), .Z(n14826) );
  CMXI2X1 U25920 ( .A0(n14826), .A1(n14820), .S(n4155), .Z(n14833) );
  CMX2X1 U25921 ( .A0(n14821), .A1(n14833), .S(n3806), .Z(n14849) );
  CMXI2X1 U25922 ( .A0(n14822), .A1(n14849), .S(n3370), .Z(N9003) );
  CMX2X1 U25923 ( .A0(N7541), .A1(N7540), .S(n3868), .Z(n14829) );
  CMXI2X1 U25924 ( .A0(n14829), .A1(n14823), .S(n4155), .Z(n14836) );
  CMX2X1 U25925 ( .A0(n14824), .A1(n14836), .S(n4305), .Z(n14852) );
  CMXI2X1 U25926 ( .A0(n14825), .A1(n14852), .S(n3370), .Z(N9004) );
  CMX2X1 U25927 ( .A0(N7540), .A1(N7539), .S(n3869), .Z(n14832) );
  CMXI2X1 U25928 ( .A0(n14832), .A1(n14826), .S(n4155), .Z(n14839) );
  CMX2X1 U25929 ( .A0(n14827), .A1(n14839), .S(n3771), .Z(n14855) );
  CMXI2X1 U25930 ( .A0(n14828), .A1(n14855), .S(n3370), .Z(N9005) );
  CMX2X1 U25931 ( .A0(N7539), .A1(N7538), .S(n3870), .Z(n14835) );
  CMXI2X1 U25932 ( .A0(n14835), .A1(n14829), .S(n4155), .Z(n14845) );
  CMX2X1 U25933 ( .A0(n14830), .A1(n14845), .S(n3772), .Z(n14858) );
  CMXI2X1 U25934 ( .A0(n14831), .A1(n14858), .S(n3370), .Z(N9006) );
  CMX2X1 U25935 ( .A0(N7538), .A1(N7537), .S(n3871), .Z(n14838) );
  CMXI2X1 U25936 ( .A0(n14838), .A1(n14832), .S(n4155), .Z(n14848) );
  CMX2X1 U25937 ( .A0(n14833), .A1(n14848), .S(n3807), .Z(n14861) );
  CMXI2X1 U25938 ( .A0(n14834), .A1(n14861), .S(n3373), .Z(N9007) );
  CMX2X1 U25939 ( .A0(N7537), .A1(N7536), .S(n3872), .Z(n14844) );
  CMXI2X1 U25940 ( .A0(n14844), .A1(n14835), .S(n4155), .Z(n14851) );
  CMX2X1 U25941 ( .A0(n14836), .A1(n14851), .S(n3808), .Z(n14864) );
  CMXI2X1 U25942 ( .A0(n14837), .A1(n14864), .S(n3373), .Z(N9008) );
  CMX2X1 U25943 ( .A0(N7536), .A1(N7535), .S(n3868), .Z(n14847) );
  CMXI2X1 U25944 ( .A0(n14847), .A1(n14838), .S(n4155), .Z(n14854) );
  CMX2X1 U25945 ( .A0(n14839), .A1(n14854), .S(n3809), .Z(n14867) );
  CMXI2X1 U25946 ( .A0(n14840), .A1(n14867), .S(n3373), .Z(N9009) );
  CMX2X1 U25947 ( .A0(N8193), .A1(N8192), .S(n3869), .Z(n14907) );
  CMXI2X1 U25948 ( .A0(n14907), .A1(n14841), .S(n4155), .Z(n14974) );
  CMX2X1 U25949 ( .A0(n14842), .A1(n14974), .S(n3810), .Z(n15111) );
  CMXI2X1 U25950 ( .A0(n14843), .A1(n15111), .S(n3373), .Z(N8352) );
  CMX2X1 U25951 ( .A0(N7535), .A1(N7534), .S(n3873), .Z(n14850) );
  CMXI2X1 U25952 ( .A0(n14850), .A1(n14844), .S(n4155), .Z(n14857) );
  CMX2X1 U25953 ( .A0(n14845), .A1(n14857), .S(n3811), .Z(n14870) );
  CMXI2X1 U25954 ( .A0(n14846), .A1(n14870), .S(n3373), .Z(N9010) );
  CMX2X1 U25955 ( .A0(N7534), .A1(N7533), .S(n3874), .Z(n14853) );
  CMXI2X1 U25956 ( .A0(n14853), .A1(n14847), .S(n4155), .Z(n14860) );
  CMX2X1 U25957 ( .A0(n14848), .A1(n14860), .S(n3812), .Z(n14873) );
  CMXI2X1 U25958 ( .A0(n14849), .A1(n14873), .S(n3373), .Z(N9011) );
  CMX2X1 U25959 ( .A0(N7533), .A1(N7532), .S(n3881), .Z(n14856) );
  CMXI2X1 U25960 ( .A0(n14856), .A1(n14850), .S(n4155), .Z(n14863) );
  CMX2X1 U25961 ( .A0(n14851), .A1(n14863), .S(n4305), .Z(n14879) );
  CMXI2X1 U25962 ( .A0(n14852), .A1(n14879), .S(n3373), .Z(N9012) );
  CMX2X1 U25963 ( .A0(N7532), .A1(N7531), .S(n3862), .Z(n14859) );
  CMXI2X1 U25964 ( .A0(n14859), .A1(n14853), .S(n4155), .Z(n14866) );
  CMX2X1 U25965 ( .A0(n14854), .A1(n14866), .S(n3771), .Z(n14882) );
  CMXI2X1 U25966 ( .A0(n14855), .A1(n14882), .S(n3372), .Z(N9013) );
  CMX2X1 U25967 ( .A0(N7531), .A1(N7530), .S(n3863), .Z(n14862) );
  CMXI2X1 U25968 ( .A0(n14862), .A1(n14856), .S(n4155), .Z(n14869) );
  CMX2X1 U25969 ( .A0(n14857), .A1(n14869), .S(n3772), .Z(n14885) );
  CMXI2X1 U25970 ( .A0(n14858), .A1(n14885), .S(n3372), .Z(N9014) );
  CMX2X1 U25971 ( .A0(N7530), .A1(N7529), .S(n3864), .Z(n14865) );
  CMXI2X1 U25972 ( .A0(n14865), .A1(n14859), .S(n4154), .Z(n14872) );
  CMX2X1 U25973 ( .A0(n14860), .A1(n14872), .S(n3773), .Z(n14888) );
  CMXI2X1 U25974 ( .A0(n14861), .A1(n14888), .S(n3372), .Z(N9015) );
  CMX2X1 U25975 ( .A0(N7529), .A1(N7528), .S(n3879), .Z(n14868) );
  CMXI2X1 U25976 ( .A0(n14868), .A1(n14862), .S(n4154), .Z(n14878) );
  CMX2X1 U25977 ( .A0(n14863), .A1(n14878), .S(n3774), .Z(n14891) );
  CMXI2X1 U25978 ( .A0(n14864), .A1(n14891), .S(n3372), .Z(N9016) );
  CMX2X1 U25979 ( .A0(N7528), .A1(N7527), .S(n3880), .Z(n14871) );
  CMXI2X1 U25980 ( .A0(n14871), .A1(n14865), .S(n4154), .Z(n14881) );
  CMX2X1 U25981 ( .A0(n14866), .A1(n14881), .S(n3775), .Z(n14894) );
  CMXI2X1 U25982 ( .A0(n14867), .A1(n14894), .S(n3372), .Z(N9017) );
  CMX2X1 U25983 ( .A0(N7527), .A1(N7526), .S(n3881), .Z(n14877) );
  CMXI2X1 U25984 ( .A0(n14877), .A1(n14868), .S(n4154), .Z(n14884) );
  CMX2X1 U25985 ( .A0(n14869), .A1(n14884), .S(n3776), .Z(n14897) );
  CMXI2X1 U25986 ( .A0(n14870), .A1(n14897), .S(n3372), .Z(N9018) );
  CMX2X1 U25987 ( .A0(N7526), .A1(N7525), .S(n3862), .Z(n14880) );
  CMXI2X1 U25988 ( .A0(n14880), .A1(n14871), .S(n4154), .Z(n14887) );
  CMX2X1 U25989 ( .A0(n14872), .A1(n14887), .S(n3777), .Z(n14900) );
  CMXI2X1 U25990 ( .A0(n14873), .A1(n14900), .S(n3372), .Z(N9019) );
  CMX2X1 U25991 ( .A0(N8192), .A1(N8191), .S(n3871), .Z(n14940) );
  CMXI2X1 U25992 ( .A0(n14940), .A1(n14874), .S(n4154), .Z(n15007) );
  CMX2X1 U25993 ( .A0(n14875), .A1(n15007), .S(n3790), .Z(n15144) );
  CMXI2X1 U25994 ( .A0(n14876), .A1(n15144), .S(n3372), .Z(N8353) );
  CMX2X1 U25995 ( .A0(N7525), .A1(N7524), .S(n3875), .Z(n14883) );
  CMXI2X1 U25996 ( .A0(n14883), .A1(n14877), .S(n4154), .Z(n14890) );
  CMX2X1 U25997 ( .A0(n14878), .A1(n14890), .S(n3791), .Z(n14903) );
  CMXI2X1 U25998 ( .A0(n14879), .A1(n14903), .S(n3372), .Z(N9020) );
  CMX2X1 U25999 ( .A0(N7524), .A1(N7523), .S(n3876), .Z(n14886) );
  CMXI2X1 U26000 ( .A0(n14886), .A1(n14880), .S(n4154), .Z(n14893) );
  CMX2X1 U26001 ( .A0(n14881), .A1(n14893), .S(n3797), .Z(n14906) );
  CMXI2X1 U26002 ( .A0(n14882), .A1(n14906), .S(n3372), .Z(N9021) );
  CMX2X1 U26003 ( .A0(N7523), .A1(N7522), .S(n3877), .Z(n14889) );
  CMXI2X1 U26004 ( .A0(n14889), .A1(n14883), .S(n4154), .Z(n14896) );
  CMX2X1 U26005 ( .A0(n14884), .A1(n14896), .S(n3774), .Z(n14912) );
  CMXI2X1 U26006 ( .A0(n14885), .A1(n14912), .S(n3375), .Z(N9022) );
  CMX2X1 U26007 ( .A0(N7522), .A1(N7521), .S(n3878), .Z(n14892) );
  CMXI2X1 U26008 ( .A0(n14892), .A1(n14886), .S(n4154), .Z(n14899) );
  CMX2X1 U26009 ( .A0(n14887), .A1(n14899), .S(n3776), .Z(n14915) );
  CMXI2X1 U26010 ( .A0(n14888), .A1(n14915), .S(n3375), .Z(N9023) );
  CMX2X1 U26011 ( .A0(N7521), .A1(N7520), .S(n3879), .Z(n14895) );
  CMXI2X1 U26012 ( .A0(n14895), .A1(n14889), .S(n4154), .Z(n14902) );
  CMX2X1 U26013 ( .A0(n14890), .A1(n14902), .S(n3777), .Z(n14918) );
  CMXI2X1 U26014 ( .A0(n14891), .A1(n14918), .S(n3375), .Z(N9024) );
  CMX2X1 U26015 ( .A0(N7520), .A1(N7519), .S(n3880), .Z(n14898) );
  CMXI2X1 U26016 ( .A0(n14898), .A1(n14892), .S(n4154), .Z(n14905) );
  CMX2X1 U26017 ( .A0(n14893), .A1(n14905), .S(n3790), .Z(n14921) );
  CMXI2X1 U26018 ( .A0(n14894), .A1(n14921), .S(n3374), .Z(N9025) );
  CMX2X1 U26019 ( .A0(N7519), .A1(N7518), .S(n3881), .Z(n14901) );
  CMXI2X1 U26020 ( .A0(n14901), .A1(n14895), .S(n4154), .Z(n14911) );
  CMX2X1 U26021 ( .A0(n14896), .A1(n14911), .S(n3791), .Z(n14924) );
  CMXI2X1 U26022 ( .A0(n14897), .A1(n14924), .S(n3374), .Z(N9026) );
  CMX2X1 U26023 ( .A0(N7518), .A1(N7517), .S(n3870), .Z(n14904) );
  CMXI2X1 U26024 ( .A0(n14904), .A1(n14898), .S(n4154), .Z(n14914) );
  CMX2X1 U26025 ( .A0(n14899), .A1(n14914), .S(n3792), .Z(n14927) );
  CMXI2X1 U26026 ( .A0(n14900), .A1(n14927), .S(n3374), .Z(N9027) );
  CMX2X1 U26027 ( .A0(N7517), .A1(N7516), .S(n3871), .Z(n14910) );
  CMXI2X1 U26028 ( .A0(n14910), .A1(n14901), .S(n4154), .Z(n14917) );
  CMX2X1 U26029 ( .A0(n14902), .A1(n14917), .S(n3793), .Z(n14930) );
  CMXI2X1 U26030 ( .A0(n14903), .A1(n14930), .S(n3374), .Z(N9028) );
  CMX2X1 U26031 ( .A0(N7516), .A1(N7515), .S(n3862), .Z(n14913) );
  CMXI2X1 U26032 ( .A0(n14913), .A1(n14904), .S(n4154), .Z(n14920) );
  CMX2X1 U26033 ( .A0(n14905), .A1(n14920), .S(n3794), .Z(n14933) );
  CMXI2X1 U26034 ( .A0(n14906), .A1(n14933), .S(n3374), .Z(N9029) );
  CMX2X1 U26035 ( .A0(N8191), .A1(N8190), .S(n3863), .Z(n14973) );
  CMXI2X1 U26036 ( .A0(n14973), .A1(n14907), .S(n4153), .Z(n15040) );
  CMX2X1 U26037 ( .A0(n14908), .A1(n15040), .S(n3795), .Z(n15177) );
  CMXI2X1 U26038 ( .A0(n14909), .A1(n15177), .S(n3374), .Z(N8354) );
  CMX2X1 U26039 ( .A0(N7515), .A1(N7514), .S(n3865), .Z(n14916) );
  CMXI2X1 U26040 ( .A0(n14916), .A1(n14910), .S(n4153), .Z(n14923) );
  CMX2X1 U26041 ( .A0(n14911), .A1(n14923), .S(n3796), .Z(n14936) );
  CMXI2X1 U26042 ( .A0(n14912), .A1(n14936), .S(n3374), .Z(N9030) );
  CMX2X1 U26043 ( .A0(N7514), .A1(N7513), .S(n3866), .Z(n14919) );
  CMXI2X1 U26044 ( .A0(n14919), .A1(n14913), .S(n4153), .Z(n14926) );
  CMX2X1 U26045 ( .A0(n14914), .A1(n14926), .S(n3797), .Z(n14939) );
  CMXI2X1 U26046 ( .A0(n14915), .A1(n14939), .S(n3374), .Z(N9031) );
  CMX2X1 U26047 ( .A0(N7513), .A1(N7512), .S(n3867), .Z(n14922) );
  CMXI2X1 U26048 ( .A0(n14922), .A1(n14916), .S(n4153), .Z(n14929) );
  CMX2X1 U26049 ( .A0(n14917), .A1(n14929), .S(n3805), .Z(n14945) );
  CMXI2X1 U26050 ( .A0(n14918), .A1(n14945), .S(n3374), .Z(N9032) );
  CMX2X1 U26051 ( .A0(N7512), .A1(N7511), .S(n3868), .Z(n14925) );
  CMXI2X1 U26052 ( .A0(n14925), .A1(n14919), .S(n4153), .Z(n14932) );
  CMX2X1 U26053 ( .A0(n14920), .A1(n14932), .S(n3806), .Z(n14948) );
  CMXI2X1 U26054 ( .A0(n14921), .A1(n14948), .S(n3374), .Z(N9033) );
  CMX2X1 U26055 ( .A0(N7511), .A1(N7510), .S(n3863), .Z(n14928) );
  CMXI2X1 U26056 ( .A0(n14928), .A1(n14922), .S(n4153), .Z(n14935) );
  CMX2X1 U26057 ( .A0(n14923), .A1(n14935), .S(n3806), .Z(n14951) );
  CMXI2X1 U26058 ( .A0(n14924), .A1(n14951), .S(n3374), .Z(N9034) );
  CMX2X1 U26059 ( .A0(N7510), .A1(N7509), .S(n3864), .Z(n14931) );
  CMXI2X1 U26060 ( .A0(n14931), .A1(n14925), .S(n4153), .Z(n14938) );
  CMX2X1 U26061 ( .A0(n14926), .A1(n14938), .S(n3791), .Z(n14954) );
  CMXI2X1 U26062 ( .A0(n14927), .A1(n14954), .S(n3373), .Z(N9035) );
  CMX2X1 U26063 ( .A0(N7509), .A1(N7508), .S(n3865), .Z(n14934) );
  CMXI2X1 U26064 ( .A0(n14934), .A1(n14928), .S(n4153), .Z(n14944) );
  CMX2X1 U26065 ( .A0(n14929), .A1(n14944), .S(n3772), .Z(n14957) );
  CMXI2X1 U26066 ( .A0(n14930), .A1(n14957), .S(n3373), .Z(N9036) );
  CMX2X1 U26067 ( .A0(N7508), .A1(N7507), .S(n3866), .Z(n14937) );
  CMXI2X1 U26068 ( .A0(n14937), .A1(n14931), .S(n4153), .Z(n14947) );
  CMX2X1 U26069 ( .A0(n14932), .A1(n14947), .S(n3773), .Z(n14960) );
  CMXI2X1 U26070 ( .A0(n14933), .A1(n14960), .S(n3373), .Z(N9037) );
  CMX2X1 U26071 ( .A0(N7507), .A1(N7506), .S(n3872), .Z(n14943) );
  CMXI2X1 U26072 ( .A0(n14943), .A1(n14934), .S(n4153), .Z(n14950) );
  CMX2X1 U26073 ( .A0(n14935), .A1(n14950), .S(n3774), .Z(n14963) );
  CMXI2X1 U26074 ( .A0(n14936), .A1(n14963), .S(n3373), .Z(N9038) );
  CMX2X1 U26075 ( .A0(N7506), .A1(N7505), .S(n3864), .Z(n14946) );
  CMXI2X1 U26076 ( .A0(n14946), .A1(n14937), .S(n4153), .Z(n14953) );
  CMX2X1 U26077 ( .A0(n14938), .A1(n14953), .S(n3775), .Z(n14966) );
  CMXI2X1 U26078 ( .A0(n14939), .A1(n14966), .S(n3376), .Z(N9039) );
  CMX2X1 U26079 ( .A0(N8190), .A1(N8189), .S(n3865), .Z(n15006) );
  CMXI2X1 U26080 ( .A0(n15006), .A1(n14940), .S(n4153), .Z(n15073) );
  CMX2X1 U26081 ( .A0(n14941), .A1(n15073), .S(n3776), .Z(n15210) );
  CMXI2X1 U26082 ( .A0(n14942), .A1(n15210), .S(n3376), .Z(N8355) );
  CMX2X1 U26083 ( .A0(N7505), .A1(N7504), .S(n3866), .Z(n14949) );
  CMXI2X1 U26084 ( .A0(n14949), .A1(n14943), .S(n4153), .Z(n14956) );
  CMX2X1 U26085 ( .A0(n14944), .A1(n14956), .S(n4306), .Z(n14969) );
  CMXI2X1 U26086 ( .A0(n14945), .A1(n14969), .S(n3376), .Z(N9040) );
  CMX2X1 U26087 ( .A0(N7504), .A1(N7503), .S(n3867), .Z(n14952) );
  CMXI2X1 U26088 ( .A0(n14952), .A1(n14946), .S(n4153), .Z(n14959) );
  CMX2X1 U26089 ( .A0(n14947), .A1(n14959), .S(n3807), .Z(n14972) );
  CMXI2X1 U26090 ( .A0(n14948), .A1(n14972), .S(n3376), .Z(N9041) );
  CMX2X1 U26091 ( .A0(N7503), .A1(N7502), .S(n3868), .Z(n14955) );
  CMXI2X1 U26092 ( .A0(n14955), .A1(n14949), .S(n4153), .Z(n14962) );
  CMX2X1 U26093 ( .A0(n14950), .A1(n14962), .S(n3808), .Z(n14978) );
  CMXI2X1 U26094 ( .A0(n14951), .A1(n14978), .S(n3376), .Z(N9042) );
  CMX2X1 U26095 ( .A0(N7502), .A1(N7501), .S(n3869), .Z(n14958) );
  CMXI2X1 U26096 ( .A0(n14958), .A1(n14952), .S(n4153), .Z(n14965) );
  CMX2X1 U26097 ( .A0(n14953), .A1(n14965), .S(n3809), .Z(n14981) );
  CMXI2X1 U26098 ( .A0(n14954), .A1(n14981), .S(n3376), .Z(N9043) );
  CMX2X1 U26099 ( .A0(N7501), .A1(N7500), .S(n3870), .Z(n14961) );
  CMXI2X1 U26100 ( .A0(n14961), .A1(n14955), .S(n4152), .Z(n14968) );
  CMX2X1 U26101 ( .A0(n14956), .A1(n14968), .S(n3810), .Z(n14984) );
  CMXI2X1 U26102 ( .A0(n14957), .A1(n14984), .S(n3376), .Z(N9044) );
  CMX2X1 U26103 ( .A0(N7500), .A1(N7499), .S(n3872), .Z(n14964) );
  CMXI2X1 U26104 ( .A0(n14964), .A1(n14958), .S(n4152), .Z(n14971) );
  CMX2X1 U26105 ( .A0(n14959), .A1(n14971), .S(n3811), .Z(n14987) );
  CMXI2X1 U26106 ( .A0(n14960), .A1(n14987), .S(n3376), .Z(N9045) );
  CMX2X1 U26107 ( .A0(N7499), .A1(N7498), .S(n3873), .Z(n14967) );
  CMXI2X1 U26108 ( .A0(n14967), .A1(n14961), .S(n4152), .Z(n14977) );
  CMX2X1 U26109 ( .A0(n14962), .A1(n14977), .S(n3812), .Z(n14990) );
  CMXI2X1 U26110 ( .A0(n14963), .A1(n14990), .S(n3376), .Z(N9046) );
  CMX2X1 U26111 ( .A0(N7498), .A1(N7497), .S(n3871), .Z(n14970) );
  CMXI2X1 U26112 ( .A0(n14970), .A1(n14964), .S(n4152), .Z(n14980) );
  CMX2X1 U26113 ( .A0(n14965), .A1(n14980), .S(n4306), .Z(n14993) );
  CMXI2X1 U26114 ( .A0(n14966), .A1(n14993), .S(n3376), .Z(N9047) );
  CMX2X1 U26115 ( .A0(N7497), .A1(N7496), .S(n3872), .Z(n14976) );
  CMXI2X1 U26116 ( .A0(n14976), .A1(n14967), .S(n4152), .Z(n14983) );
  CMX2X1 U26117 ( .A0(n14968), .A1(n14983), .S(n3771), .Z(n14996) );
  CMXI2X1 U26118 ( .A0(n14969), .A1(n14996), .S(n3375), .Z(N9048) );
  CMX2X1 U26119 ( .A0(N7496), .A1(N7495), .S(n3869), .Z(n14979) );
  CMXI2X1 U26120 ( .A0(n14979), .A1(n14970), .S(n4152), .Z(n14986) );
  CMX2X1 U26121 ( .A0(n14971), .A1(n14986), .S(n3772), .Z(n14999) );
  CMXI2X1 U26122 ( .A0(n14972), .A1(n14999), .S(n3375), .Z(N9049) );
  CMX2X1 U26123 ( .A0(N8189), .A1(N8188), .S(n3870), .Z(n15039) );
  CMXI2X1 U26124 ( .A0(n15039), .A1(n14973), .S(n4152), .Z(n15110) );
  CMX2X1 U26125 ( .A0(n14974), .A1(n15110), .S(n3773), .Z(n15243) );
  CMXI2X1 U26126 ( .A0(n14975), .A1(n15243), .S(n3375), .Z(N8356) );
  CMX2X1 U26127 ( .A0(N7495), .A1(N7494), .S(n3871), .Z(n14982) );
  CMXI2X1 U26128 ( .A0(n14982), .A1(n14976), .S(n4152), .Z(n14989) );
  CMX2X1 U26129 ( .A0(n14977), .A1(n14989), .S(n3774), .Z(n15002) );
  CMXI2X1 U26130 ( .A0(n14978), .A1(n15002), .S(n3375), .Z(N9050) );
  CMX2X1 U26131 ( .A0(N7494), .A1(N7493), .S(n3872), .Z(n14985) );
  CMXI2X1 U26132 ( .A0(n14985), .A1(n14979), .S(n4152), .Z(n14992) );
  CMX2X1 U26133 ( .A0(n14980), .A1(n14992), .S(n3775), .Z(n15005) );
  CMXI2X1 U26134 ( .A0(n14981), .A1(n15005), .S(n3375), .Z(N9051) );
  CMX2X1 U26135 ( .A0(N7493), .A1(N7492), .S(n3867), .Z(n14988) );
  CMXI2X1 U26136 ( .A0(n14988), .A1(n14982), .S(n4152), .Z(n14995) );
  CMX2X1 U26137 ( .A0(n14983), .A1(n14995), .S(n3776), .Z(n15011) );
  CMXI2X1 U26138 ( .A0(n14984), .A1(n15011), .S(n3375), .Z(N9052) );
  CMX2X1 U26139 ( .A0(N7492), .A1(N7491), .S(n3868), .Z(n14991) );
  CMXI2X1 U26140 ( .A0(n14991), .A1(n14985), .S(n4152), .Z(n14998) );
  CMX2X1 U26141 ( .A0(n14986), .A1(n14998), .S(n3777), .Z(n15014) );
  CMXI2X1 U26142 ( .A0(n14987), .A1(n15014), .S(n3375), .Z(N9053) );
  CMX2X1 U26143 ( .A0(N7491), .A1(N7490), .S(n3869), .Z(n14994) );
  CMXI2X1 U26144 ( .A0(n14994), .A1(n14988), .S(n4152), .Z(n15001) );
  CMX2X1 U26145 ( .A0(n14989), .A1(n15001), .S(n3790), .Z(n15017) );
  CMXI2X1 U26146 ( .A0(n14990), .A1(n15017), .S(n3375), .Z(N9054) );
  CMX2X1 U26147 ( .A0(N7490), .A1(N7489), .S(n3870), .Z(n14997) );
  CMXI2X1 U26148 ( .A0(n14997), .A1(n14991), .S(n4152), .Z(n15004) );
  CMX2X1 U26149 ( .A0(n14992), .A1(n15004), .S(n3791), .Z(n15020) );
  CMXI2X1 U26150 ( .A0(n14993), .A1(n15020), .S(n3378), .Z(N9055) );
  CMX2X1 U26151 ( .A0(N7489), .A1(N7488), .S(n3873), .Z(n15000) );
  CMXI2X1 U26152 ( .A0(n15000), .A1(n14994), .S(n4152), .Z(n15010) );
  CMX2X1 U26153 ( .A0(n14995), .A1(n15010), .S(n3807), .Z(n15023) );
  CMXI2X1 U26154 ( .A0(n14996), .A1(n15023), .S(n3378), .Z(N9056) );
  CMX2X1 U26155 ( .A0(N7488), .A1(N7487), .S(n3873), .Z(n15003) );
  CMXI2X1 U26156 ( .A0(n15003), .A1(n14997), .S(n4152), .Z(n15013) );
  CMX2X1 U26157 ( .A0(n14998), .A1(n15013), .S(n3792), .Z(n15026) );
  CMXI2X1 U26158 ( .A0(n14999), .A1(n15026), .S(n3378), .Z(N9057) );
  CMX2X1 U26159 ( .A0(N7487), .A1(N7486), .S(n3874), .Z(n15009) );
  CMXI2X1 U26160 ( .A0(n15009), .A1(n15000), .S(n4152), .Z(n15016) );
  CMX2X1 U26161 ( .A0(n15001), .A1(n15016), .S(n3777), .Z(n15029) );
  CMXI2X1 U26162 ( .A0(n15002), .A1(n15029), .S(n3378), .Z(N9058) );
  CMX2X1 U26163 ( .A0(N7486), .A1(N7485), .S(n3875), .Z(n15012) );
  CMXI2X1 U26164 ( .A0(n15012), .A1(n15003), .S(n4151), .Z(n15019) );
  CMX2X1 U26165 ( .A0(n15004), .A1(n15019), .S(n3790), .Z(n15032) );
  CMXI2X1 U26166 ( .A0(n15005), .A1(n15032), .S(n3378), .Z(N9059) );
  CMX2X1 U26167 ( .A0(N8188), .A1(N8187), .S(n3876), .Z(n15072) );
  CMXI2X1 U26168 ( .A0(n15072), .A1(n15006), .S(n4151), .Z(n15143) );
  CMX2X1 U26169 ( .A0(n15007), .A1(n15143), .S(n3791), .Z(n15276) );
  CMXI2X1 U26170 ( .A0(n15008), .A1(n15276), .S(n3378), .Z(N8357) );
  CMX2X1 U26171 ( .A0(N7485), .A1(N7484), .S(n3877), .Z(n15015) );
  CMXI2X1 U26172 ( .A0(n15015), .A1(n15009), .S(n4151), .Z(n15022) );
  CMX2X1 U26173 ( .A0(n15010), .A1(n15022), .S(n3792), .Z(n15035) );
  CMXI2X1 U26174 ( .A0(n15011), .A1(n15035), .S(n3377), .Z(N9060) );
  CMX2X1 U26175 ( .A0(N7484), .A1(N7483), .S(n3878), .Z(n15018) );
  CMXI2X1 U26176 ( .A0(n15018), .A1(n15012), .S(n4151), .Z(n15025) );
  CMX2X1 U26177 ( .A0(n15013), .A1(n15025), .S(n3793), .Z(n15038) );
  CMXI2X1 U26178 ( .A0(n15014), .A1(n15038), .S(n3377), .Z(N9061) );
  CMX2X1 U26179 ( .A0(N7483), .A1(N7482), .S(n3879), .Z(n15021) );
  CMXI2X1 U26180 ( .A0(n15021), .A1(n15015), .S(n4151), .Z(n15028) );
  CMX2X1 U26181 ( .A0(n15016), .A1(n15028), .S(n3771), .Z(n15044) );
  CMXI2X1 U26182 ( .A0(n15017), .A1(n15044), .S(n3377), .Z(N9062) );
  CMX2X1 U26183 ( .A0(N7482), .A1(N7481), .S(n3874), .Z(n15024) );
  CMXI2X1 U26184 ( .A0(n15024), .A1(n15018), .S(n4151), .Z(n15031) );
  CMX2X1 U26185 ( .A0(n15019), .A1(n15031), .S(n3792), .Z(n15047) );
  CMXI2X1 U26186 ( .A0(n15020), .A1(n15047), .S(n3377), .Z(N9063) );
  CMX2X1 U26187 ( .A0(N7481), .A1(N7480), .S(n3875), .Z(n15027) );
  CMXI2X1 U26188 ( .A0(n15027), .A1(n15021), .S(n4151), .Z(n15034) );
  CMX2X1 U26189 ( .A0(n15022), .A1(n15034), .S(n3793), .Z(n15050) );
  CMXI2X1 U26190 ( .A0(n15023), .A1(n15050), .S(n3377), .Z(N9064) );
  CMX2X1 U26191 ( .A0(N7480), .A1(N7479), .S(n3880), .Z(n15030) );
  CMXI2X1 U26192 ( .A0(n15030), .A1(n15024), .S(n4151), .Z(n15037) );
  CMX2X1 U26193 ( .A0(n15025), .A1(n15037), .S(n3794), .Z(n15053) );
  CMXI2X1 U26194 ( .A0(n15026), .A1(n15053), .S(n3377), .Z(N9065) );
  CMX2X1 U26195 ( .A0(N7479), .A1(N7478), .S(n3881), .Z(n15033) );
  CMXI2X1 U26196 ( .A0(n15033), .A1(n15027), .S(n4151), .Z(n15043) );
  CMX2X1 U26197 ( .A0(n15028), .A1(n15043), .S(n3795), .Z(n15056) );
  CMXI2X1 U26198 ( .A0(n15029), .A1(n15056), .S(n3377), .Z(N9066) );
  CMX2X1 U26199 ( .A0(N7478), .A1(N7477), .S(n3873), .Z(n15036) );
  CMXI2X1 U26200 ( .A0(n15036), .A1(n15030), .S(n4151), .Z(n15046) );
  CMX2X1 U26201 ( .A0(n15031), .A1(n15046), .S(n3796), .Z(n15059) );
  CMXI2X1 U26202 ( .A0(n15032), .A1(n15059), .S(n3377), .Z(N9067) );
  CMX2X1 U26203 ( .A0(N7477), .A1(N7476), .S(n3874), .Z(n15042) );
  CMXI2X1 U26204 ( .A0(n15042), .A1(n15033), .S(n4151), .Z(n15049) );
  CMX2X1 U26205 ( .A0(n15034), .A1(n15049), .S(n3797), .Z(n15062) );
  CMXI2X1 U26206 ( .A0(n15035), .A1(n15062), .S(n3377), .Z(N9068) );
  CMX2X1 U26207 ( .A0(N7476), .A1(N7475), .S(n3875), .Z(n15045) );
  CMXI2X1 U26208 ( .A0(n15045), .A1(n15036), .S(n4151), .Z(n15052) );
  CMX2X1 U26209 ( .A0(n15037), .A1(n15052), .S(n3805), .Z(n15065) );
  CMXI2X1 U26210 ( .A0(n15038), .A1(n15065), .S(n3377), .Z(N9069) );
  CMX2X1 U26211 ( .A0(N8187), .A1(N8186), .S(n3876), .Z(n15109) );
  CMXI2X1 U26212 ( .A0(n15109), .A1(n15039), .S(n4151), .Z(n15176) );
  CMX2X1 U26213 ( .A0(n15040), .A1(n15176), .S(n3806), .Z(n15310) );
  CMXI2X1 U26214 ( .A0(n15041), .A1(n15310), .S(n3377), .Z(N8358) );
  CMX2X1 U26215 ( .A0(N7475), .A1(N7474), .S(n3871), .Z(n15048) );
  CMXI2X1 U26216 ( .A0(n15048), .A1(n15042), .S(n4151), .Z(n15055) );
  CMX2X1 U26217 ( .A0(n15043), .A1(n15055), .S(n3807), .Z(n15068) );
  CMXI2X1 U26218 ( .A0(n15044), .A1(n15068), .S(n3376), .Z(N9070) );
  CMX2X1 U26219 ( .A0(N7474), .A1(N7473), .S(n3872), .Z(n15051) );
  CMXI2X1 U26220 ( .A0(n15051), .A1(n15045), .S(n4151), .Z(n15058) );
  CMX2X1 U26221 ( .A0(n15046), .A1(n15058), .S(n3808), .Z(n15071) );
  CMXI2X1 U26222 ( .A0(n15047), .A1(n15071), .S(n3380), .Z(N9071) );
  CMX2X1 U26223 ( .A0(N7473), .A1(N7472), .S(n3873), .Z(n15054) );
  CMXI2X1 U26224 ( .A0(n15054), .A1(n15048), .S(n4151), .Z(n15061) );
  CMX2X1 U26225 ( .A0(n15049), .A1(n15061), .S(n3809), .Z(n15081) );
  CMXI2X1 U26226 ( .A0(n15050), .A1(n15081), .S(n3380), .Z(N9072) );
  CMX2X1 U26227 ( .A0(N7472), .A1(N7471), .S(n3874), .Z(n15057) );
  CMXI2X1 U26228 ( .A0(n15057), .A1(n15051), .S(n4150), .Z(n15064) );
  CMX2X1 U26229 ( .A0(n15052), .A1(n15064), .S(n3810), .Z(n15084) );
  CMXI2X1 U26230 ( .A0(n15053), .A1(n15084), .S(n3379), .Z(N9073) );
  CMX2X1 U26231 ( .A0(N7471), .A1(N7470), .S(n3874), .Z(n15060) );
  CMXI2X1 U26232 ( .A0(n15060), .A1(n15054), .S(n4150), .Z(n15067) );
  CMX2X1 U26233 ( .A0(n15055), .A1(n15067), .S(n3811), .Z(n15087) );
  CMXI2X1 U26234 ( .A0(n15056), .A1(n15087), .S(n3379), .Z(N9074) );
  CMX2X1 U26235 ( .A0(N7470), .A1(N7469), .S(n3862), .Z(n15063) );
  CMXI2X1 U26236 ( .A0(n15063), .A1(n15057), .S(n4150), .Z(n15070) );
  CMX2X1 U26237 ( .A0(n15058), .A1(n15070), .S(n3812), .Z(n15090) );
  CMXI2X1 U26238 ( .A0(n15059), .A1(n15090), .S(n3379), .Z(N9075) );
  CMX2X1 U26239 ( .A0(N7469), .A1(N7468), .S(n3863), .Z(n15066) );
  CMXI2X1 U26240 ( .A0(n15066), .A1(n15060), .S(n4150), .Z(n15080) );
  CMX2X1 U26241 ( .A0(n15061), .A1(n15080), .S(n4305), .Z(n15093) );
  CMXI2X1 U26242 ( .A0(n15062), .A1(n15093), .S(n3379), .Z(N9076) );
  CMX2X1 U26243 ( .A0(N7468), .A1(N7467), .S(n3864), .Z(n15069) );
  CMXI2X1 U26244 ( .A0(n15069), .A1(n15063), .S(n4150), .Z(n15083) );
  CMX2X1 U26245 ( .A0(n15064), .A1(n15083), .S(n3771), .Z(n15096) );
  CMXI2X1 U26246 ( .A0(n15065), .A1(n15096), .S(n3379), .Z(N9077) );
  CMX2X1 U26247 ( .A0(N7467), .A1(N7466), .S(n3865), .Z(n15079) );
  CMXI2X1 U26248 ( .A0(n15079), .A1(n15066), .S(n4150), .Z(n15086) );
  CMX2X1 U26249 ( .A0(n15067), .A1(n15086), .S(n3808), .Z(n15099) );
  CMXI2X1 U26250 ( .A0(n15068), .A1(n15099), .S(n3379), .Z(N9078) );
  CMX2X1 U26251 ( .A0(N7466), .A1(N7465), .S(n3866), .Z(n15082) );
  CMXI2X1 U26252 ( .A0(n15082), .A1(n15069), .S(n4150), .Z(n15089) );
  CMX2X1 U26253 ( .A0(n15070), .A1(n15089), .S(n3793), .Z(n15102) );
  CMXI2X1 U26254 ( .A0(n15071), .A1(n15102), .S(n3379), .Z(N9079) );
  CMX2X1 U26255 ( .A0(N8186), .A1(N8185), .S(n3865), .Z(n15142) );
  CMXI2X1 U26256 ( .A0(n15142), .A1(n15072), .S(n4150), .Z(n15209) );
  CMX2X1 U26257 ( .A0(n15073), .A1(n15209), .S(n3794), .Z(n15344) );
  CMXI2X1 U26258 ( .A0(n15074), .A1(n15344), .S(n3379), .Z(N8359) );
  CMXI2X1 U26259 ( .A0(n15078), .A1(n15077), .S(n3379), .Z(N8287) );
  CMX2X1 U26260 ( .A0(N7465), .A1(N7464), .S(n3876), .Z(n15085) );
  CMXI2X1 U26261 ( .A0(n15085), .A1(n15079), .S(n4150), .Z(n15092) );
  CMX2X1 U26262 ( .A0(n15080), .A1(n15092), .S(n3795), .Z(n15105) );
  CMXI2X1 U26263 ( .A0(n15081), .A1(n15105), .S(n3379), .Z(N9080) );
  CMX2X1 U26264 ( .A0(N7464), .A1(N7463), .S(n3877), .Z(n15088) );
  CMXI2X1 U26265 ( .A0(n15088), .A1(n15082), .S(n4150), .Z(n15095) );
  CMX2X1 U26266 ( .A0(n15083), .A1(n15095), .S(n3796), .Z(n15108) );
  CMXI2X1 U26267 ( .A0(n15084), .A1(n15108), .S(n3379), .Z(N9081) );
  CMX2X1 U26268 ( .A0(N7463), .A1(N7462), .S(n3869), .Z(n15091) );
  CMXI2X1 U26269 ( .A0(n15091), .A1(n15085), .S(n4150), .Z(n15098) );
  CMX2X1 U26270 ( .A0(n15086), .A1(n15098), .S(n3797), .Z(n15114) );
  CMXI2X1 U26271 ( .A0(n15087), .A1(n15114), .S(n3378), .Z(N9082) );
  CMX2X1 U26272 ( .A0(N7462), .A1(N7461), .S(n3870), .Z(n15094) );
  CMXI2X1 U26273 ( .A0(n15094), .A1(n15088), .S(n4150), .Z(n15101) );
  CMX2X1 U26274 ( .A0(n15089), .A1(n15101), .S(n3805), .Z(n15117) );
  CMXI2X1 U26275 ( .A0(n15090), .A1(n15117), .S(n3378), .Z(N9083) );
  CMX2X1 U26276 ( .A0(N7461), .A1(N7460), .S(n3871), .Z(n15097) );
  CMXI2X1 U26277 ( .A0(n15097), .A1(n15091), .S(n4150), .Z(n15104) );
  CMX2X1 U26278 ( .A0(n15092), .A1(n15104), .S(n3772), .Z(n15120) );
  CMXI2X1 U26279 ( .A0(n15093), .A1(n15120), .S(n3378), .Z(N9084) );
  CMX2X1 U26280 ( .A0(N7460), .A1(N7459), .S(n3872), .Z(n15100) );
  CMXI2X1 U26281 ( .A0(n15100), .A1(n15094), .S(n4150), .Z(n15107) );
  CMX2X1 U26282 ( .A0(n15095), .A1(n15107), .S(n3772), .Z(n15123) );
  CMXI2X1 U26283 ( .A0(n15096), .A1(n15123), .S(n3378), .Z(N9085) );
  CMX2X1 U26284 ( .A0(N7459), .A1(N7458), .S(n3867), .Z(n15103) );
  CMXI2X1 U26285 ( .A0(n15103), .A1(n15097), .S(n4150), .Z(n15113) );
  CMX2X1 U26286 ( .A0(n15098), .A1(n15113), .S(n3773), .Z(n15126) );
  CMXI2X1 U26287 ( .A0(n15099), .A1(n15126), .S(n3378), .Z(N9086) );
  CMX2X1 U26288 ( .A0(N7458), .A1(N7457), .S(n3868), .Z(n15106) );
  CMXI2X1 U26289 ( .A0(n15106), .A1(n15100), .S(n4150), .Z(n15116) );
  CMX2X1 U26290 ( .A0(n15101), .A1(n15116), .S(n3774), .Z(n15129) );
  CMXI2X1 U26291 ( .A0(n15102), .A1(n15129), .S(n3479), .Z(N9087) );
  CMX2X1 U26292 ( .A0(N7457), .A1(N7456), .S(n3869), .Z(n15112) );
  CMXI2X1 U26293 ( .A0(n15112), .A1(n15103), .S(n4149), .Z(n15119) );
  CMX2X1 U26294 ( .A0(n15104), .A1(n15119), .S(n3775), .Z(n15132) );
  CMXI2X1 U26295 ( .A0(n15105), .A1(n15132), .S(n3515), .Z(N9088) );
  CMX2X1 U26296 ( .A0(N7456), .A1(N7455), .S(n3870), .Z(n15115) );
  CMXI2X1 U26297 ( .A0(n15115), .A1(n15106), .S(n4149), .Z(n15122) );
  CMX2X1 U26298 ( .A0(n15107), .A1(n15122), .S(n3776), .Z(n15135) );
  CMXI2X1 U26299 ( .A0(n15108), .A1(n15135), .S(n3482), .Z(N9089) );
  CMX2X1 U26300 ( .A0(N8185), .A1(N8184), .S(n3878), .Z(n15175) );
  CMXI2X1 U26301 ( .A0(n15175), .A1(n15109), .S(n4149), .Z(n15242) );
  CMX2X1 U26302 ( .A0(n15110), .A1(n15242), .S(n3777), .Z(n15377) );
  CMXI2X1 U26303 ( .A0(n15111), .A1(n15377), .S(n3360), .Z(N8360) );
  CMX2X1 U26304 ( .A0(N7455), .A1(N7454), .S(n3878), .Z(n15118) );
  CMXI2X1 U26305 ( .A0(n15118), .A1(n15112), .S(n4149), .Z(n15125) );
  CMX2X1 U26306 ( .A0(n15113), .A1(n15125), .S(n3790), .Z(n15138) );
  CMXI2X1 U26307 ( .A0(n15114), .A1(n15138), .S(n3517), .Z(N9090) );
  CMX2X1 U26308 ( .A0(N7454), .A1(N7453), .S(n3879), .Z(n15121) );
  CMXI2X1 U26309 ( .A0(n15121), .A1(n15115), .S(n4149), .Z(n15128) );
  CMX2X1 U26310 ( .A0(n15116), .A1(n15128), .S(n3793), .Z(n15141) );
  CMXI2X1 U26311 ( .A0(n15117), .A1(n15141), .S(n3516), .Z(N9091) );
  CMX2X1 U26312 ( .A0(N7453), .A1(N7452), .S(n3880), .Z(n15124) );
  CMXI2X1 U26313 ( .A0(n15124), .A1(n15118), .S(n4149), .Z(n15131) );
  CMX2X1 U26314 ( .A0(n15119), .A1(n15131), .S(n3772), .Z(n15147) );
  CMXI2X1 U26315 ( .A0(n15120), .A1(n15147), .S(n3498), .Z(N9092) );
  CMX2X1 U26316 ( .A0(N7452), .A1(N7451), .S(n3881), .Z(n15127) );
  CMXI2X1 U26317 ( .A0(n15127), .A1(n15121), .S(n4149), .Z(n15134) );
  CMX2X1 U26318 ( .A0(n15122), .A1(n15134), .S(n3773), .Z(n15150) );
  CMXI2X1 U26319 ( .A0(n15123), .A1(n15150), .S(n3497), .Z(N9093) );
  CMX2X1 U26320 ( .A0(N7451), .A1(N7450), .S(n3862), .Z(n15130) );
  CMXI2X1 U26321 ( .A0(n15130), .A1(n15124), .S(n4149), .Z(n15137) );
  CMX2X1 U26322 ( .A0(n15125), .A1(n15137), .S(n3774), .Z(n15153) );
  CMXI2X1 U26323 ( .A0(n15126), .A1(n15153), .S(n3380), .Z(N9094) );
  CMX2X1 U26324 ( .A0(N7450), .A1(N7449), .S(n3863), .Z(n15133) );
  CMXI2X1 U26325 ( .A0(n15133), .A1(n15127), .S(n4149), .Z(n15140) );
  CMX2X1 U26326 ( .A0(n15128), .A1(n15140), .S(n3775), .Z(n15156) );
  CMXI2X1 U26327 ( .A0(n15129), .A1(n15156), .S(n3380), .Z(N9095) );
  CMX2X1 U26328 ( .A0(N7449), .A1(N7448), .S(n3864), .Z(n15136) );
  CMXI2X1 U26329 ( .A0(n15136), .A1(n15130), .S(n4149), .Z(n15146) );
  CMX2X1 U26330 ( .A0(n15131), .A1(n15146), .S(n3776), .Z(n15159) );
  CMXI2X1 U26331 ( .A0(n15132), .A1(n15159), .S(n3380), .Z(N9096) );
  CMX2X1 U26332 ( .A0(N7448), .A1(N7447), .S(n3864), .Z(n15139) );
  CMXI2X1 U26333 ( .A0(n15139), .A1(n15133), .S(n4149), .Z(n15149) );
  CMX2X1 U26334 ( .A0(n15134), .A1(n15149), .S(n3777), .Z(n15162) );
  CMXI2X1 U26335 ( .A0(n15135), .A1(n15162), .S(n3380), .Z(N9097) );
  CMX2X1 U26336 ( .A0(N7447), .A1(N7446), .S(n3865), .Z(n15145) );
  CMXI2X1 U26337 ( .A0(n15145), .A1(n15136), .S(n4149), .Z(n15152) );
  CMX2X1 U26338 ( .A0(n15137), .A1(n15152), .S(n3790), .Z(n15165) );
  CMXI2X1 U26339 ( .A0(n15138), .A1(n15165), .S(n3380), .Z(N9098) );
  CMX2X1 U26340 ( .A0(N7446), .A1(N7445), .S(n3865), .Z(n15148) );
  CMXI2X1 U26341 ( .A0(n15148), .A1(n15139), .S(n4149), .Z(n15155) );
  CMX2X1 U26342 ( .A0(n15140), .A1(n15155), .S(n3791), .Z(n15168) );
  CMXI2X1 U26343 ( .A0(n15141), .A1(n15168), .S(n3380), .Z(N9099) );
  CMX2X1 U26344 ( .A0(N8184), .A1(N8183), .S(n3866), .Z(n15208) );
  CMXI2X1 U26345 ( .A0(n15208), .A1(n15142), .S(n4149), .Z(n15275) );
  CMX2X1 U26346 ( .A0(n15143), .A1(n15275), .S(n3791), .Z(n15410) );
  CMXI2X1 U26347 ( .A0(n15144), .A1(n15410), .S(n3380), .Z(N8361) );
  CMX2X1 U26348 ( .A0(N7445), .A1(N7444), .S(n3873), .Z(n15151) );
  CMXI2X1 U26349 ( .A0(n15151), .A1(n15145), .S(n4149), .Z(n15158) );
  CMX2X1 U26350 ( .A0(n15146), .A1(n15158), .S(n3771), .Z(n15171) );
  CMXI2X1 U26351 ( .A0(n15147), .A1(n15171), .S(n3380), .Z(N9100) );
  CMX2X1 U26352 ( .A0(N7444), .A1(N7443), .S(n3874), .Z(n15154) );
  CMXI2X1 U26353 ( .A0(n15154), .A1(n15148), .S(n4149), .Z(n15161) );
  CMX2X1 U26354 ( .A0(n15149), .A1(n15161), .S(n3792), .Z(n15174) );
  CMXI2X1 U26355 ( .A0(n15150), .A1(n15174), .S(n3380), .Z(N9101) );
  CMX2X1 U26356 ( .A0(N7443), .A1(N7442), .S(n3875), .Z(n15157) );
  CMXI2X1 U26357 ( .A0(n15157), .A1(n15151), .S(n4148), .Z(n15164) );
  CMX2X1 U26358 ( .A0(n15152), .A1(n15164), .S(n3793), .Z(n15180) );
  CMXI2X1 U26359 ( .A0(n15153), .A1(n15180), .S(n3394), .Z(N9102) );
  CMX2X1 U26360 ( .A0(N7442), .A1(N7441), .S(n3876), .Z(n15160) );
  CMXI2X1 U26361 ( .A0(n15160), .A1(n15154), .S(n4148), .Z(n15167) );
  CMX2X1 U26362 ( .A0(n15155), .A1(n15167), .S(n3794), .Z(n15183) );
  CMXI2X1 U26363 ( .A0(n15156), .A1(n15183), .S(n3486), .Z(N9103) );
  CMX2X1 U26364 ( .A0(N7441), .A1(N7440), .S(n3871), .Z(n15163) );
  CMXI2X1 U26365 ( .A0(n15163), .A1(n15157), .S(n4148), .Z(n15170) );
  CMX2X1 U26366 ( .A0(n15158), .A1(n15170), .S(n3795), .Z(n15186) );
  CMXI2X1 U26367 ( .A0(n15159), .A1(n15186), .S(n3485), .Z(N9104) );
  CMX2X1 U26368 ( .A0(N7440), .A1(N7439), .S(n3872), .Z(n15166) );
  CMXI2X1 U26369 ( .A0(n15166), .A1(n15160), .S(n4148), .Z(n15173) );
  CMX2X1 U26370 ( .A0(n15161), .A1(n15173), .S(n3796), .Z(n15189) );
  CMXI2X1 U26371 ( .A0(n15162), .A1(n15189), .S(n3484), .Z(N9105) );
  CMX2X1 U26372 ( .A0(N7439), .A1(N7438), .S(n3873), .Z(n15169) );
  CMXI2X1 U26373 ( .A0(n15169), .A1(n15163), .S(n4148), .Z(n15179) );
  CMX2X1 U26374 ( .A0(n15164), .A1(n15179), .S(n3805), .Z(n15192) );
  CMXI2X1 U26375 ( .A0(n15165), .A1(n15192), .S(n3483), .Z(N9106) );
  CMX2X1 U26376 ( .A0(N7438), .A1(N7437), .S(n3874), .Z(n15172) );
  CMXI2X1 U26377 ( .A0(n15172), .A1(n15166), .S(n4148), .Z(n15182) );
  CMX2X1 U26378 ( .A0(n15167), .A1(n15182), .S(n3792), .Z(n15195) );
  CMXI2X1 U26379 ( .A0(n15168), .A1(n15195), .S(n3380), .Z(N9107) );
  CMX2X1 U26380 ( .A0(N7437), .A1(N7436), .S(n3879), .Z(n15178) );
  CMXI2X1 U26381 ( .A0(n15178), .A1(n15169), .S(n4148), .Z(n15185) );
  CMX2X1 U26382 ( .A0(n15170), .A1(n15185), .S(n3807), .Z(n15198) );
  CMXI2X1 U26383 ( .A0(n15171), .A1(n15198), .S(n3387), .Z(N9108) );
  CMX2X1 U26384 ( .A0(N7436), .A1(N7435), .S(n3867), .Z(n15181) );
  CMXI2X1 U26385 ( .A0(n15181), .A1(n15172), .S(n4148), .Z(n15188) );
  CMX2X1 U26386 ( .A0(n15173), .A1(n15188), .S(n3808), .Z(n15201) );
  CMXI2X1 U26387 ( .A0(n15174), .A1(n15201), .S(n3350), .Z(N9109) );
  CMX2X1 U26388 ( .A0(N8183), .A1(N8182), .S(n3868), .Z(n15241) );
  CMXI2X1 U26389 ( .A0(n15241), .A1(n15175), .S(n4148), .Z(n15309) );
  CMX2X1 U26390 ( .A0(n15176), .A1(n15309), .S(n3809), .Z(n15445) );
  CMXI2X1 U26391 ( .A0(n15177), .A1(n15445), .S(n3367), .Z(N8362) );
  CMX2X1 U26392 ( .A0(N7435), .A1(N7434), .S(n3869), .Z(n15184) );
  CMXI2X1 U26393 ( .A0(n15184), .A1(n15178), .S(n4148), .Z(n15191) );
  CMX2X1 U26394 ( .A0(n15179), .A1(n15191), .S(n3810), .Z(n15204) );
  CMXI2X1 U26395 ( .A0(n15180), .A1(n15204), .S(n3349), .Z(N9110) );
  CMX2X1 U26396 ( .A0(N7434), .A1(N7433), .S(n3870), .Z(n15187) );
  CMXI2X1 U26397 ( .A0(n15187), .A1(n15181), .S(n4148), .Z(n15194) );
  CMX2X1 U26398 ( .A0(n15182), .A1(n15194), .S(n3811), .Z(n15207) );
  CMXI2X1 U26399 ( .A0(n15183), .A1(n15207), .S(n3348), .Z(N9111) );
  CMX2X1 U26400 ( .A0(N7433), .A1(N7432), .S(n3871), .Z(n15190) );
  CMXI2X1 U26401 ( .A0(n15190), .A1(n15184), .S(n4148), .Z(n15197) );
  CMX2X1 U26402 ( .A0(n15185), .A1(n15197), .S(n3812), .Z(n15213) );
  CMXI2X1 U26403 ( .A0(n15186), .A1(n15213), .S(n3493), .Z(N9112) );
  CMX2X1 U26404 ( .A0(N7432), .A1(N7431), .S(n3872), .Z(n15193) );
  CMXI2X1 U26405 ( .A0(n15193), .A1(n15187), .S(n4148), .Z(n15200) );
  CMX2X1 U26406 ( .A0(n15188), .A1(n15200), .S(n4305), .Z(n15216) );
  CMXI2X1 U26407 ( .A0(n15189), .A1(n15216), .S(n3351), .Z(N9113) );
  CMX2X1 U26408 ( .A0(N7431), .A1(N7430), .S(n3873), .Z(n15196) );
  CMXI2X1 U26409 ( .A0(n15196), .A1(n15190), .S(n4148), .Z(n15203) );
  CMX2X1 U26410 ( .A0(n15191), .A1(n15203), .S(n3771), .Z(n15219) );
  CMXI2X1 U26411 ( .A0(n15192), .A1(n15219), .S(n3345), .Z(N9114) );
  CMX2X1 U26412 ( .A0(N7430), .A1(N7429), .S(n3866), .Z(n15199) );
  CMXI2X1 U26413 ( .A0(n15199), .A1(n15193), .S(n4148), .Z(n15206) );
  CMX2X1 U26414 ( .A0(n15194), .A1(n15206), .S(n3771), .Z(n15222) );
  CMXI2X1 U26415 ( .A0(n15195), .A1(n15222), .S(n3344), .Z(N9115) );
  CMX2X1 U26416 ( .A0(N7429), .A1(N7428), .S(n3867), .Z(n15202) );
  CMXI2X1 U26417 ( .A0(n15202), .A1(n15196), .S(n4148), .Z(n15212) );
  CMX2X1 U26418 ( .A0(n15197), .A1(n15212), .S(n3806), .Z(n15225) );
  CMXI2X1 U26419 ( .A0(n15198), .A1(n15225), .S(n3343), .Z(N9116) );
  CMX2X1 U26420 ( .A0(N7428), .A1(N7427), .S(n3874), .Z(n15205) );
  CMXI2X1 U26421 ( .A0(n15205), .A1(n15199), .S(n4147), .Z(n15215) );
  CMX2X1 U26422 ( .A0(n15200), .A1(n15215), .S(n3807), .Z(n15228) );
  CMXI2X1 U26423 ( .A0(n15201), .A1(n15228), .S(n3342), .Z(N9117) );
  CMX2X1 U26424 ( .A0(N7427), .A1(N7426), .S(n3875), .Z(n15211) );
  CMXI2X1 U26425 ( .A0(n15211), .A1(n15202), .S(n4147), .Z(n15218) );
  CMX2X1 U26426 ( .A0(n15203), .A1(n15218), .S(n3808), .Z(n15231) );
  CMXI2X1 U26427 ( .A0(n15204), .A1(n15231), .S(n3341), .Z(N9118) );
  CMX2X1 U26428 ( .A0(N7426), .A1(N7425), .S(n3877), .Z(n15214) );
  CMXI2X1 U26429 ( .A0(n15214), .A1(n15205), .S(n4147), .Z(n15221) );
  CMX2X1 U26430 ( .A0(n15206), .A1(n15221), .S(n3809), .Z(n15234) );
  CMXI2X1 U26431 ( .A0(n15207), .A1(n15234), .S(n3340), .Z(N9119) );
  CMX2X1 U26432 ( .A0(N8182), .A1(N8181), .S(n3878), .Z(n15274) );
  CMXI2X1 U26433 ( .A0(n15274), .A1(n15208), .S(n4147), .Z(n15343) );
  CMX2X1 U26434 ( .A0(n15209), .A1(n15343), .S(n3810), .Z(n15478) );
  CMXI2X1 U26435 ( .A0(n15210), .A1(n15478), .S(n3339), .Z(N8363) );
  CMX2X1 U26436 ( .A0(N7425), .A1(N7424), .S(n3879), .Z(n15217) );
  CMXI2X1 U26437 ( .A0(n15217), .A1(n15211), .S(n4147), .Z(n15224) );
  CMX2X1 U26438 ( .A0(n15212), .A1(n15224), .S(n3811), .Z(n15237) );
  CMXI2X1 U26439 ( .A0(n15213), .A1(n15237), .S(n3338), .Z(N9120) );
  CMX2X1 U26440 ( .A0(N7424), .A1(N7423), .S(n3880), .Z(n15220) );
  CMXI2X1 U26441 ( .A0(n15220), .A1(n15214), .S(n4147), .Z(n15227) );
  CMX2X1 U26442 ( .A0(n15215), .A1(n15227), .S(n3790), .Z(n15240) );
  CMXI2X1 U26443 ( .A0(n15216), .A1(n15240), .S(n3337), .Z(N9121) );
  CMX2X1 U26444 ( .A0(N7423), .A1(N7422), .S(n3875), .Z(n15223) );
  CMXI2X1 U26445 ( .A0(n15223), .A1(n15217), .S(n4147), .Z(n15230) );
  CMX2X1 U26446 ( .A0(n15218), .A1(n15230), .S(n3772), .Z(n15246) );
  CMXI2X1 U26447 ( .A0(n15219), .A1(n15246), .S(n3372), .Z(N9122) );
  CMX2X1 U26448 ( .A0(N7422), .A1(N7421), .S(n3876), .Z(n15226) );
  CMXI2X1 U26449 ( .A0(n15226), .A1(n15220), .S(n4147), .Z(n15233) );
  CMX2X1 U26450 ( .A0(n15221), .A1(n15233), .S(n3773), .Z(n15249) );
  CMXI2X1 U26451 ( .A0(n15222), .A1(n15249), .S(n3370), .Z(N9123) );
  CMX2X1 U26452 ( .A0(N7421), .A1(N7420), .S(n3877), .Z(n15229) );
  CMXI2X1 U26453 ( .A0(n15229), .A1(n15223), .S(n4147), .Z(n15236) );
  CMX2X1 U26454 ( .A0(n15224), .A1(n15236), .S(n3774), .Z(n15252) );
  CMXI2X1 U26455 ( .A0(n15225), .A1(n15252), .S(n3369), .Z(N9124) );
  CMX2X1 U26456 ( .A0(N7420), .A1(N7419), .S(n3878), .Z(n15232) );
  CMXI2X1 U26457 ( .A0(n15232), .A1(n15226), .S(n4147), .Z(n15239) );
  CMX2X1 U26458 ( .A0(n15227), .A1(n15239), .S(n3775), .Z(n15255) );
  CMXI2X1 U26459 ( .A0(n15228), .A1(n15255), .S(n3378), .Z(N9125) );
  CMX2X1 U26460 ( .A0(N7419), .A1(N7418), .S(n3880), .Z(n15235) );
  CMXI2X1 U26461 ( .A0(n15235), .A1(n15229), .S(n4147), .Z(n15245) );
  CMX2X1 U26462 ( .A0(n15230), .A1(n15245), .S(n3776), .Z(n15258) );
  CMXI2X1 U26463 ( .A0(n15231), .A1(n15258), .S(n3377), .Z(N9126) );
  CMX2X1 U26464 ( .A0(N7418), .A1(N7417), .S(n3876), .Z(n15238) );
  CMXI2X1 U26465 ( .A0(n15238), .A1(n15232), .S(n4147), .Z(n15248) );
  CMX2X1 U26466 ( .A0(n15233), .A1(n15248), .S(n3777), .Z(n15261) );
  CMXI2X1 U26467 ( .A0(n15234), .A1(n15261), .S(n3376), .Z(N9127) );
  CMX2X1 U26468 ( .A0(N7417), .A1(N7416), .S(n3877), .Z(n15244) );
  CMXI2X1 U26469 ( .A0(n15244), .A1(n15235), .S(n4147), .Z(n15251) );
  CMX2X1 U26470 ( .A0(n15236), .A1(n15251), .S(n3790), .Z(n15264) );
  CMXI2X1 U26471 ( .A0(n15237), .A1(n15264), .S(n3375), .Z(N9128) );
  CMX2X1 U26472 ( .A0(N7416), .A1(N7415), .S(n3878), .Z(n15247) );
  CMXI2X1 U26473 ( .A0(n15247), .A1(n15238), .S(n4147), .Z(n15254) );
  CMX2X1 U26474 ( .A0(n15239), .A1(n15254), .S(n3791), .Z(n15267) );
  CMXI2X1 U26475 ( .A0(n15240), .A1(n15267), .S(n3374), .Z(N9129) );
  CMX2X1 U26476 ( .A0(N8181), .A1(N8180), .S(n3879), .Z(n15307) );
  CMXI2X1 U26477 ( .A0(n15307), .A1(n15241), .S(n4147), .Z(n15376) );
  CMX2X1 U26478 ( .A0(n15242), .A1(n15376), .S(n3792), .Z(n15510) );
  CMXI2X1 U26479 ( .A0(n15243), .A1(n15510), .S(n3373), .Z(N8364) );
  CMX2X1 U26480 ( .A0(N7415), .A1(N7414), .S(n3880), .Z(n15250) );
  CMXI2X1 U26481 ( .A0(n15250), .A1(n15244), .S(n4147), .Z(n15257) );
  CMX2X1 U26482 ( .A0(n15245), .A1(n15257), .S(n3793), .Z(n15270) );
  CMXI2X1 U26483 ( .A0(n15246), .A1(n15270), .S(n3347), .Z(N9130) );
  CMX2X1 U26484 ( .A0(N7414), .A1(N7413), .S(n3881), .Z(n15253) );
  CMXI2X1 U26485 ( .A0(n15253), .A1(n15247), .S(n4146), .Z(n15260) );
  CMX2X1 U26486 ( .A0(n15248), .A1(n15260), .S(n3794), .Z(n15273) );
  CMXI2X1 U26487 ( .A0(n15249), .A1(n15273), .S(n3346), .Z(N9131) );
  CMX2X1 U26488 ( .A0(N7413), .A1(N7412), .S(n3862), .Z(n15256) );
  CMXI2X1 U26489 ( .A0(n15256), .A1(n15250), .S(n4146), .Z(n15263) );
  CMX2X1 U26490 ( .A0(n15251), .A1(n15263), .S(n3795), .Z(n15279) );
  CMXI2X1 U26491 ( .A0(n15252), .A1(n15279), .S(n3336), .Z(N9132) );
  CMX2X1 U26492 ( .A0(N7412), .A1(N7411), .S(n3868), .Z(n15259) );
  CMXI2X1 U26493 ( .A0(n15259), .A1(n15253), .S(n4146), .Z(n15266) );
  CMX2X1 U26494 ( .A0(n15254), .A1(n15266), .S(n3796), .Z(n15282) );
  CMXI2X1 U26495 ( .A0(n15255), .A1(n15282), .S(n3332), .Z(N9133) );
  CMX2X1 U26496 ( .A0(N7411), .A1(N7410), .S(n3869), .Z(n15262) );
  CMXI2X1 U26497 ( .A0(n15262), .A1(n15256), .S(n4146), .Z(n15269) );
  CMX2X1 U26498 ( .A0(n15257), .A1(n15269), .S(n3797), .Z(n15285) );
  CMXI2X1 U26499 ( .A0(n15258), .A1(n15285), .S(n3518), .Z(N9134) );
  CMX2X1 U26500 ( .A0(N7410), .A1(N7409), .S(n3863), .Z(n15265) );
  CMXI2X1 U26501 ( .A0(n15265), .A1(n15259), .S(n4146), .Z(n15272) );
  CMX2X1 U26502 ( .A0(n15260), .A1(n15272), .S(n3805), .Z(n15288) );
  CMXI2X1 U26503 ( .A0(n15261), .A1(n15288), .S(n3364), .Z(N9135) );
  CMX2X1 U26504 ( .A0(N7409), .A1(N7408), .S(n3864), .Z(n15268) );
  CMXI2X1 U26505 ( .A0(n15268), .A1(n15262), .S(n4146), .Z(n15278) );
  CMX2X1 U26506 ( .A0(n15263), .A1(n15278), .S(n3806), .Z(n15291) );
  CMXI2X1 U26507 ( .A0(n15264), .A1(n15291), .S(n3363), .Z(N9136) );
  CMX2X1 U26508 ( .A0(N7408), .A1(N7407), .S(n3881), .Z(n15271) );
  CMXI2X1 U26509 ( .A0(n15271), .A1(n15265), .S(n4146), .Z(n15281) );
  CMX2X1 U26510 ( .A0(n15266), .A1(n15281), .S(n3772), .Z(n15294) );
  CMXI2X1 U26511 ( .A0(n15267), .A1(n15294), .S(n3362), .Z(N9137) );
  CMX2X1 U26512 ( .A0(N7407), .A1(N7406), .S(n3862), .Z(n15277) );
  CMXI2X1 U26513 ( .A0(n15277), .A1(n15268), .S(n4146), .Z(n15284) );
  CMX2X1 U26514 ( .A0(n15269), .A1(n15284), .S(n3807), .Z(n15297) );
  CMXI2X1 U26515 ( .A0(n15270), .A1(n15297), .S(n3361), .Z(N9138) );
  CMX2X1 U26516 ( .A0(N7406), .A1(N7405), .S(n3863), .Z(n15280) );
  CMXI2X1 U26517 ( .A0(n15280), .A1(n15271), .S(n4146), .Z(n15287) );
  CMX2X1 U26518 ( .A0(n15272), .A1(n15287), .S(n3812), .Z(n15300) );
  CMXI2X1 U26519 ( .A0(n15273), .A1(n15300), .S(n3366), .Z(N9139) );
  CMX2X1 U26520 ( .A0(N8180), .A1(N8179), .S(n3864), .Z(n15341) );
  CMXI2X1 U26521 ( .A0(n15341), .A1(n15274), .S(n4146), .Z(n15409) );
  CMX2X1 U26522 ( .A0(n15275), .A1(n15409), .S(n4306), .Z(n15542) );
  CMXI2X1 U26523 ( .A0(n15276), .A1(n15542), .S(n3368), .Z(N8365) );
  CMX2X1 U26524 ( .A0(N7405), .A1(N7404), .S(n3879), .Z(n15283) );
  CMXI2X1 U26525 ( .A0(n15283), .A1(n15277), .S(n4146), .Z(n15290) );
  CMX2X1 U26526 ( .A0(n15278), .A1(n15290), .S(n3771), .Z(n15303) );
  CMXI2X1 U26527 ( .A0(n15279), .A1(n15303), .S(n3365), .Z(N9140) );
  CMX2X1 U26528 ( .A0(N7404), .A1(N7403), .S(n3880), .Z(n15286) );
  CMXI2X1 U26529 ( .A0(n15286), .A1(n15280), .S(n4146), .Z(n15293) );
  CMX2X1 U26530 ( .A0(n15281), .A1(n15293), .S(n3772), .Z(n15306) );
  CMXI2X1 U26531 ( .A0(n15282), .A1(n15306), .S(n3382), .Z(N9141) );
  CMX2X1 U26532 ( .A0(N7403), .A1(N7402), .S(n3881), .Z(n15289) );
  CMXI2X1 U26533 ( .A0(n15289), .A1(n15283), .S(n4146), .Z(n15296) );
  CMX2X1 U26534 ( .A0(n15284), .A1(n15296), .S(n3773), .Z(n15313) );
  CMXI2X1 U26535 ( .A0(n15285), .A1(n15313), .S(n3382), .Z(N9142) );
  CMX2X1 U26536 ( .A0(N7402), .A1(N7401), .S(n3862), .Z(n15292) );
  CMXI2X1 U26537 ( .A0(n15292), .A1(n15286), .S(n4146), .Z(n15299) );
  CMX2X1 U26538 ( .A0(n15287), .A1(n15299), .S(n3791), .Z(n15316) );
  CMXI2X1 U26539 ( .A0(n15288), .A1(n15316), .S(n3382), .Z(N9143) );
  CMX2X1 U26540 ( .A0(N7401), .A1(N7400), .S(n3881), .Z(n15295) );
  CMXI2X1 U26541 ( .A0(n15295), .A1(n15289), .S(n4146), .Z(n15302) );
  CMX2X1 U26542 ( .A0(n15290), .A1(n15302), .S(n3807), .Z(n15319) );
  CMXI2X1 U26543 ( .A0(n15291), .A1(n15319), .S(n3382), .Z(N9144) );
  CMX2X1 U26544 ( .A0(N7400), .A1(N7399), .S(n3865), .Z(n15298) );
  CMXI2X1 U26545 ( .A0(n15298), .A1(n15292), .S(n4146), .Z(n15305) );
  CMX2X1 U26546 ( .A0(n15293), .A1(n15305), .S(n3808), .Z(n15322) );
  CMXI2X1 U26547 ( .A0(n15294), .A1(n15322), .S(n3382), .Z(N9145) );
  CMX2X1 U26548 ( .A0(N7399), .A1(N7398), .S(n3866), .Z(n15301) );
  CMXI2X1 U26549 ( .A0(n15301), .A1(n15295), .S(n4145), .Z(n15312) );
  CMX2X1 U26550 ( .A0(n15296), .A1(n15312), .S(n3809), .Z(n15325) );
  CMXI2X1 U26551 ( .A0(n15297), .A1(n15325), .S(n3382), .Z(N9146) );
  CMX2X1 U26552 ( .A0(N7398), .A1(N7397), .S(n3867), .Z(n15304) );
  CMXI2X1 U26553 ( .A0(n15304), .A1(n15298), .S(n4145), .Z(n15315) );
  CMX2X1 U26554 ( .A0(n15299), .A1(n15315), .S(n3810), .Z(n15328) );
  CMXI2X1 U26555 ( .A0(n15300), .A1(n15328), .S(n3382), .Z(N9147) );
  CMX2X1 U26556 ( .A0(N7397), .A1(N7396), .S(n3868), .Z(n15311) );
  CMXI2X1 U26557 ( .A0(n15311), .A1(n15301), .S(n4145), .Z(n15318) );
  CMX2X1 U26558 ( .A0(n15302), .A1(n15318), .S(n3811), .Z(n15331) );
  CMXI2X1 U26559 ( .A0(n15303), .A1(n15331), .S(n3381), .Z(N9148) );
  CMX2X1 U26560 ( .A0(N7396), .A1(N7395), .S(n3869), .Z(n15314) );
  CMXI2X1 U26561 ( .A0(n15314), .A1(n15304), .S(n4145), .Z(n15321) );
  CMX2X1 U26562 ( .A0(n15305), .A1(n15321), .S(n3812), .Z(n15334) );
  CMXI2X1 U26563 ( .A0(n15306), .A1(n15334), .S(n3381), .Z(N9149) );
  CMXI2X1 U26564 ( .A0(n15308), .A1(n15307), .S(n4145), .Z(n15444) );
  CMX2X1 U26565 ( .A0(n15309), .A1(n15444), .S(n4306), .Z(n15574) );
  CMXI2X1 U26566 ( .A0(n15310), .A1(n15574), .S(n3381), .Z(N8366) );
  CMX2X1 U26567 ( .A0(N7395), .A1(N7394), .S(n3870), .Z(n15317) );
  CMXI2X1 U26568 ( .A0(n15317), .A1(n15311), .S(n4145), .Z(n15324) );
  CMX2X1 U26569 ( .A0(n15312), .A1(n15324), .S(n3771), .Z(n15337) );
  CMXI2X1 U26570 ( .A0(n15313), .A1(n15337), .S(n3381), .Z(N9150) );
  CMX2X1 U26571 ( .A0(N7394), .A1(N7393), .S(n3871), .Z(n15320) );
  CMXI2X1 U26572 ( .A0(n15320), .A1(n15314), .S(n4145), .Z(n15327) );
  CMX2X1 U26573 ( .A0(n15315), .A1(n15327), .S(n3772), .Z(n15340) );
  CMXI2X1 U26574 ( .A0(n15316), .A1(n15340), .S(n3381), .Z(N9151) );
  CMX2X1 U26575 ( .A0(N7393), .A1(N7392), .S(n3870), .Z(n15323) );
  CMXI2X1 U26576 ( .A0(n15323), .A1(n15317), .S(n4145), .Z(n15330) );
  CMX2X1 U26577 ( .A0(n15318), .A1(n15330), .S(n3773), .Z(n15347) );
  CMXI2X1 U26578 ( .A0(n15319), .A1(n15347), .S(n3381), .Z(N9152) );
  CMX2X1 U26579 ( .A0(N7392), .A1(N7391), .S(n3871), .Z(n15326) );
  CMXI2X1 U26580 ( .A0(n15326), .A1(n15320), .S(n4145), .Z(n15333) );
  CMX2X1 U26581 ( .A0(n15321), .A1(n15333), .S(n3774), .Z(n15350) );
  CMXI2X1 U26582 ( .A0(n15322), .A1(n15350), .S(n3381), .Z(N9153) );
  CMX2X1 U26583 ( .A0(N7391), .A1(N7390), .S(n3872), .Z(n15329) );
  CMXI2X1 U26584 ( .A0(n15329), .A1(n15323), .S(n4145), .Z(n15336) );
  CMX2X1 U26585 ( .A0(n15324), .A1(n15336), .S(n3775), .Z(n15353) );
  CMXI2X1 U26586 ( .A0(n15325), .A1(n15353), .S(n3381), .Z(N9154) );
  CMX2X1 U26587 ( .A0(N7390), .A1(N7389), .S(n3873), .Z(n15332) );
  CMXI2X1 U26588 ( .A0(n15332), .A1(n15326), .S(n4145), .Z(n15339) );
  CMX2X1 U26589 ( .A0(n15327), .A1(n15339), .S(n3776), .Z(n15356) );
  CMXI2X1 U26590 ( .A0(n15328), .A1(n15356), .S(n3381), .Z(N9155) );
  CMX2X1 U26591 ( .A0(N7389), .A1(N7388), .S(n3865), .Z(n15335) );
  CMXI2X1 U26592 ( .A0(n15335), .A1(n15329), .S(n4145), .Z(n15346) );
  CMX2X1 U26593 ( .A0(n15330), .A1(n15346), .S(n3777), .Z(n15359) );
  CMXI2X1 U26594 ( .A0(n15331), .A1(n15359), .S(n3381), .Z(N9156) );
  CMX2X1 U26595 ( .A0(N7388), .A1(N7387), .S(n3866), .Z(n15338) );
  CMXI2X1 U26596 ( .A0(n15338), .A1(n15332), .S(n4145), .Z(n15349) );
  CMX2X1 U26597 ( .A0(n15333), .A1(n15349), .S(n3790), .Z(n15362) );
  CMXI2X1 U26598 ( .A0(n15334), .A1(n15362), .S(n3381), .Z(N9157) );
  CMX2X1 U26599 ( .A0(N7387), .A1(N7386), .S(n3867), .Z(n15345) );
  CMXI2X1 U26600 ( .A0(n15345), .A1(n15335), .S(n4145), .Z(n15352) );
  CMX2X1 U26601 ( .A0(n15336), .A1(n15352), .S(n3791), .Z(n15365) );
  CMXI2X1 U26602 ( .A0(n15337), .A1(n15365), .S(n3384), .Z(N9158) );
  CMX2X1 U26603 ( .A0(N7386), .A1(N7385), .S(n3868), .Z(n15348) );
  CMXI2X1 U26604 ( .A0(n15348), .A1(n15338), .S(n4145), .Z(n15355) );
  CMX2X1 U26605 ( .A0(n15339), .A1(n15355), .S(n3773), .Z(n15368) );
  CMXI2X1 U26606 ( .A0(n15340), .A1(n15368), .S(n3384), .Z(N9159) );
  CMXI2X1 U26607 ( .A0(n15342), .A1(n15341), .S(n4145), .Z(n15477) );
  CMX2X1 U26608 ( .A0(n15343), .A1(n15477), .S(n3808), .Z(n15606) );
  CMXI2X1 U26609 ( .A0(n15344), .A1(n15606), .S(n3384), .Z(N8367) );
  CMX2X1 U26610 ( .A0(N7385), .A1(N7384), .S(n3863), .Z(n15351) );
  CMXI2X1 U26611 ( .A0(n15351), .A1(n15345), .S(n4144), .Z(n15358) );
  CMX2X1 U26612 ( .A0(n15346), .A1(n15358), .S(n3774), .Z(n15371) );
  CMXI2X1 U26613 ( .A0(n15347), .A1(n15371), .S(n3383), .Z(N9160) );
  CMX2X1 U26614 ( .A0(N7384), .A1(N7383), .S(n3864), .Z(n15354) );
  CMXI2X1 U26615 ( .A0(n15354), .A1(n15348), .S(n4144), .Z(n15361) );
  CMX2X1 U26616 ( .A0(n15349), .A1(n15361), .S(n3775), .Z(n15374) );
  CMXI2X1 U26617 ( .A0(n15350), .A1(n15374), .S(n3383), .Z(N9161) );
  CMX2X1 U26618 ( .A0(N7383), .A1(N7382), .S(n3865), .Z(n15357) );
  CMXI2X1 U26619 ( .A0(n15357), .A1(n15351), .S(n4144), .Z(n15364) );
  CMX2X1 U26620 ( .A0(n15352), .A1(n15364), .S(n3776), .Z(n15380) );
  CMXI2X1 U26621 ( .A0(n15353), .A1(n15380), .S(n3383), .Z(N9162) );
  CMX2X1 U26622 ( .A0(N7382), .A1(N7381), .S(n3866), .Z(n15360) );
  CMXI2X1 U26623 ( .A0(n15360), .A1(n15354), .S(n4144), .Z(n15367) );
  CMX2X1 U26624 ( .A0(n15355), .A1(n15367), .S(n3777), .Z(n15383) );
  CMXI2X1 U26625 ( .A0(n15356), .A1(n15383), .S(n3383), .Z(N9163) );
  CMX2X1 U26626 ( .A0(N7381), .A1(N7380), .S(n3862), .Z(n15363) );
  CMXI2X1 U26627 ( .A0(n15363), .A1(n15357), .S(n4144), .Z(n15370) );
  CMX2X1 U26628 ( .A0(n15358), .A1(n15370), .S(n3790), .Z(n15386) );
  CMXI2X1 U26629 ( .A0(n15359), .A1(n15386), .S(n3383), .Z(N9164) );
  CMX2X1 U26630 ( .A0(N7380), .A1(N7379), .S(n3874), .Z(n15366) );
  CMXI2X1 U26631 ( .A0(n15366), .A1(n15360), .S(n4144), .Z(n15373) );
  CMX2X1 U26632 ( .A0(n15361), .A1(n15373), .S(n3792), .Z(n15389) );
  CMXI2X1 U26633 ( .A0(n15362), .A1(n15389), .S(n3383), .Z(N9165) );
  CMX2X1 U26634 ( .A0(N7379), .A1(N7378), .S(n3875), .Z(n15369) );
  CMXI2X1 U26635 ( .A0(n15369), .A1(n15363), .S(n4144), .Z(n15379) );
  CMX2X1 U26636 ( .A0(n15364), .A1(n15379), .S(n3792), .Z(n15392) );
  CMXI2X1 U26637 ( .A0(n15365), .A1(n15392), .S(n3383), .Z(N9166) );
  CMX2X1 U26638 ( .A0(N7378), .A1(N7377), .S(n3876), .Z(n15372) );
  CMXI2X1 U26639 ( .A0(n15372), .A1(n15366), .S(n4144), .Z(n15382) );
  CMX2X1 U26640 ( .A0(n15367), .A1(n15382), .S(n3793), .Z(n15395) );
  CMXI2X1 U26641 ( .A0(n15368), .A1(n15395), .S(n3383), .Z(N9167) );
  CMX2X1 U26642 ( .A0(N7377), .A1(N7376), .S(n3877), .Z(n15378) );
  CMXI2X1 U26643 ( .A0(n15378), .A1(n15369), .S(n4144), .Z(n15385) );
  CMX2X1 U26644 ( .A0(n15370), .A1(n15385), .S(n3794), .Z(n15398) );
  CMXI2X1 U26645 ( .A0(n15371), .A1(n15398), .S(n3383), .Z(N9168) );
  CMX2X1 U26646 ( .A0(N7376), .A1(N7375), .S(n3879), .Z(n15381) );
  CMXI2X1 U26647 ( .A0(n15381), .A1(n15372), .S(n4144), .Z(n15388) );
  CMX2X1 U26648 ( .A0(n15373), .A1(n15388), .S(n3795), .Z(n15401) );
  CMXI2X1 U26649 ( .A0(n15374), .A1(n15401), .S(n3383), .Z(N9169) );
  CMX2X1 U26650 ( .A0(n15376), .A1(n15375), .S(n3796), .Z(n15638) );
  CMXI2X1 U26651 ( .A0(n15377), .A1(n15638), .S(n3383), .Z(N8368) );
  CMX2X1 U26652 ( .A0(N7375), .A1(N7374), .S(n3880), .Z(n15384) );
  CMXI2X1 U26653 ( .A0(n15384), .A1(n15378), .S(n4144), .Z(n15391) );
  CMX2X1 U26654 ( .A0(n15379), .A1(n15391), .S(n3797), .Z(n15404) );
  CMXI2X1 U26655 ( .A0(n15380), .A1(n15404), .S(n3382), .Z(N9170) );
  CMX2X1 U26656 ( .A0(N7374), .A1(N7373), .S(n3872), .Z(n15387) );
  CMXI2X1 U26657 ( .A0(n15387), .A1(n15381), .S(n4144), .Z(n15394) );
  CMX2X1 U26658 ( .A0(n15382), .A1(n15394), .S(n3805), .Z(n15407) );
  CMXI2X1 U26659 ( .A0(n15383), .A1(n15407), .S(n3382), .Z(N9171) );
  CMX2X1 U26660 ( .A0(N7373), .A1(N7372), .S(n3873), .Z(n15390) );
  CMXI2X1 U26661 ( .A0(n15390), .A1(n15384), .S(n4144), .Z(n15397) );
  CMX2X1 U26662 ( .A0(n15385), .A1(n15397), .S(n3806), .Z(n15415) );
  CMXI2X1 U26663 ( .A0(n15386), .A1(n15415), .S(n3382), .Z(N9172) );
  CMX2X1 U26664 ( .A0(N7372), .A1(N7371), .S(n3865), .Z(n15393) );
  CMXI2X1 U26665 ( .A0(n15393), .A1(n15387), .S(n4144), .Z(n15400) );
  CMX2X1 U26666 ( .A0(n15388), .A1(n15400), .S(n3807), .Z(n15418) );
  CMXI2X1 U26667 ( .A0(n15389), .A1(n15418), .S(n3382), .Z(N9173) );
  CMX2X1 U26668 ( .A0(N7371), .A1(N7370), .S(n3866), .Z(n15396) );
  CMXI2X1 U26669 ( .A0(n15396), .A1(n15390), .S(n4144), .Z(n15403) );
  CMX2X1 U26670 ( .A0(n15391), .A1(n15403), .S(n3808), .Z(n15421) );
  CMXI2X1 U26671 ( .A0(n15392), .A1(n15421), .S(n3385), .Z(N9174) );
  CMX2X1 U26672 ( .A0(N7370), .A1(N7369), .S(n3864), .Z(n15399) );
  CMXI2X1 U26673 ( .A0(n15399), .A1(n15393), .S(n4144), .Z(n15406) );
  CMX2X1 U26674 ( .A0(n15394), .A1(n15406), .S(n3809), .Z(n15424) );
  CMXI2X1 U26675 ( .A0(n15395), .A1(n15424), .S(n3385), .Z(N9175) );
  CMX2X1 U26676 ( .A0(N7369), .A1(N7368), .S(n3865), .Z(n15402) );
  CMXI2X1 U26677 ( .A0(n15402), .A1(n15396), .S(n4143), .Z(n15414) );
  CMX2X1 U26678 ( .A0(n15397), .A1(n15414), .S(n3810), .Z(n15427) );
  CMXI2X1 U26679 ( .A0(n15398), .A1(n15427), .S(n3385), .Z(N9176) );
  CMX2X1 U26680 ( .A0(N7368), .A1(N7367), .S(n3866), .Z(n15405) );
  CMXI2X1 U26681 ( .A0(n15405), .A1(n15399), .S(n4143), .Z(n15417) );
  CMX2X1 U26682 ( .A0(n15400), .A1(n15417), .S(n3811), .Z(n15430) );
  CMXI2X1 U26683 ( .A0(n15401), .A1(n15430), .S(n3385), .Z(N9177) );
  CMX2X1 U26684 ( .A0(N7367), .A1(N7366), .S(n3867), .Z(n15413) );
  CMXI2X1 U26685 ( .A0(n15413), .A1(n15402), .S(n4143), .Z(n15420) );
  CMX2X1 U26686 ( .A0(n15403), .A1(n15420), .S(n4305), .Z(n15433) );
  CMXI2X1 U26687 ( .A0(n15404), .A1(n15433), .S(n3385), .Z(N9178) );
  CMX2X1 U26688 ( .A0(N7366), .A1(N7365), .S(n3868), .Z(n15416) );
  CMXI2X1 U26689 ( .A0(n15416), .A1(n15405), .S(n4143), .Z(n15423) );
  CMX2X1 U26690 ( .A0(n15406), .A1(n15423), .S(n3771), .Z(n15436) );
  CMXI2X1 U26691 ( .A0(n15407), .A1(n15436), .S(n3385), .Z(N9179) );
  CMX2X1 U26692 ( .A0(n15409), .A1(n15408), .S(n3774), .Z(n15670) );
  CMXI2X1 U26693 ( .A0(n15410), .A1(n15670), .S(n3385), .Z(N8369) );
  CMXI2X1 U26694 ( .A0(n15412), .A1(n15411), .S(n3385), .Z(N8288) );
  CMX2X1 U26695 ( .A0(N7365), .A1(N7364), .S(n3869), .Z(n15419) );
  CMXI2X1 U26696 ( .A0(n15419), .A1(n15413), .S(n4143), .Z(n15426) );
  CMX2X1 U26697 ( .A0(n15414), .A1(n15426), .S(n3809), .Z(n15439) );
  CMXI2X1 U26698 ( .A0(n15415), .A1(n15439), .S(n3385), .Z(N9180) );
  CMX2X1 U26699 ( .A0(N7364), .A1(N7363), .S(n3870), .Z(n15422) );
  CMXI2X1 U26700 ( .A0(n15422), .A1(n15416), .S(n4143), .Z(n15429) );
  CMX2X1 U26701 ( .A0(n15417), .A1(n15429), .S(n3791), .Z(n15442) );
  CMXI2X1 U26702 ( .A0(n15418), .A1(n15442), .S(n3385), .Z(N9181) );
  CMX2X1 U26703 ( .A0(N7363), .A1(N7362), .S(n3871), .Z(n15425) );
  CMXI2X1 U26704 ( .A0(n15425), .A1(n15419), .S(n4143), .Z(n15432) );
  CMX2X1 U26705 ( .A0(n15420), .A1(n15432), .S(n3792), .Z(n15448) );
  CMXI2X1 U26706 ( .A0(n15421), .A1(n15448), .S(n3384), .Z(N9182) );
  CMX2X1 U26707 ( .A0(N7362), .A1(N7361), .S(n3872), .Z(n15428) );
  CMXI2X1 U26708 ( .A0(n15428), .A1(n15422), .S(n4143), .Z(n15435) );
  CMX2X1 U26709 ( .A0(n15423), .A1(n15435), .S(n3793), .Z(n15451) );
  CMXI2X1 U26710 ( .A0(n15424), .A1(n15451), .S(n3384), .Z(N9183) );
  CMX2X1 U26711 ( .A0(N7361), .A1(N7360), .S(n3871), .Z(n15431) );
  CMXI2X1 U26712 ( .A0(n15431), .A1(n15425), .S(n4143), .Z(n15438) );
  CMX2X1 U26713 ( .A0(n15426), .A1(n15438), .S(n3794), .Z(n15454) );
  CMXI2X1 U26714 ( .A0(n15427), .A1(n15454), .S(n3384), .Z(N9184) );
  CMX2X1 U26715 ( .A0(N7360), .A1(N7359), .S(n3872), .Z(n15434) );
  CMXI2X1 U26716 ( .A0(n15434), .A1(n15428), .S(n4143), .Z(n15441) );
  CMX2X1 U26717 ( .A0(n15429), .A1(n15441), .S(n3795), .Z(n15457) );
  CMXI2X1 U26718 ( .A0(n15430), .A1(n15457), .S(n3384), .Z(N9185) );
  CMX2X1 U26719 ( .A0(N7359), .A1(N7358), .S(n3873), .Z(n15437) );
  CMXI2X1 U26720 ( .A0(n15437), .A1(n15431), .S(n4143), .Z(n15447) );
  CMX2X1 U26721 ( .A0(n15432), .A1(n15447), .S(n3793), .Z(n15460) );
  CMXI2X1 U26722 ( .A0(n15433), .A1(n15460), .S(n3384), .Z(N9186) );
  CMX2X1 U26723 ( .A0(N7358), .A1(N7357), .S(n3874), .Z(n15440) );
  CMXI2X1 U26724 ( .A0(n15440), .A1(n15434), .S(n4143), .Z(n15450) );
  CMX2X1 U26725 ( .A0(n15435), .A1(n15450), .S(n3772), .Z(n15463) );
  CMXI2X1 U26726 ( .A0(n15436), .A1(n15463), .S(n3384), .Z(N9187) );
  CMX2X1 U26727 ( .A0(N7357), .A1(N7356), .S(n3875), .Z(n15446) );
  CMXI2X1 U26728 ( .A0(n15446), .A1(n15437), .S(n4143), .Z(n15453) );
  CMX2X1 U26729 ( .A0(n15438), .A1(n15453), .S(n3773), .Z(n15466) );
  CMXI2X1 U26730 ( .A0(n15439), .A1(n15466), .S(n3384), .Z(N9188) );
  CMX2X1 U26731 ( .A0(N7356), .A1(N7355), .S(n3876), .Z(n15449) );
  CMXI2X1 U26732 ( .A0(n15449), .A1(n15440), .S(n4143), .Z(n15456) );
  CMX2X1 U26733 ( .A0(n15441), .A1(n15456), .S(n3774), .Z(n15469) );
  CMXI2X1 U26734 ( .A0(n15442), .A1(n15469), .S(n3384), .Z(N9189) );
  CMX2X1 U26735 ( .A0(n15444), .A1(n15443), .S(n3775), .Z(n15704) );
  CMXI2X1 U26736 ( .A0(n15445), .A1(n15704), .S(n3387), .Z(N8370) );
  CMX2X1 U26737 ( .A0(N7355), .A1(N7354), .S(n3866), .Z(n15452) );
  CMXI2X1 U26738 ( .A0(n15452), .A1(n15446), .S(n4143), .Z(n15459) );
  CMX2X1 U26739 ( .A0(n15447), .A1(n15459), .S(n3776), .Z(n15472) );
  CMXI2X1 U26740 ( .A0(n15448), .A1(n15472), .S(n3387), .Z(N9190) );
  CMX2X1 U26741 ( .A0(N7354), .A1(N7353), .S(n3867), .Z(n15455) );
  CMXI2X1 U26742 ( .A0(n15455), .A1(n15449), .S(n4143), .Z(n15462) );
  CMX2X1 U26743 ( .A0(n15450), .A1(n15462), .S(n3777), .Z(n15475) );
  CMXI2X1 U26744 ( .A0(n15451), .A1(n15475), .S(n3387), .Z(N9191) );
  CMX2X1 U26745 ( .A0(N7353), .A1(N7352), .S(n3868), .Z(n15458) );
  CMXI2X1 U26746 ( .A0(n15458), .A1(n15452), .S(n4142), .Z(n15465) );
  CMX2X1 U26747 ( .A0(n15453), .A1(n15465), .S(n3790), .Z(n15481) );
  CMXI2X1 U26748 ( .A0(n15454), .A1(n15481), .S(n3387), .Z(N9192) );
  CMX2X1 U26749 ( .A0(N7352), .A1(N7351), .S(n3869), .Z(n15461) );
  CMXI2X1 U26750 ( .A0(n15461), .A1(n15455), .S(n4142), .Z(n15468) );
  CMX2X1 U26751 ( .A0(n15456), .A1(n15468), .S(n3791), .Z(n15484) );
  CMXI2X1 U26752 ( .A0(n15457), .A1(n15484), .S(n3387), .Z(N9193) );
  CMX2X1 U26753 ( .A0(N7351), .A1(N7350), .S(n3867), .Z(n15464) );
  CMXI2X1 U26754 ( .A0(n15464), .A1(n15458), .S(n4142), .Z(n15471) );
  CMX2X1 U26755 ( .A0(n15459), .A1(n15471), .S(n3792), .Z(n15487) );
  CMXI2X1 U26756 ( .A0(n15460), .A1(n15487), .S(n3387), .Z(N9194) );
  CMX2X1 U26757 ( .A0(N7350), .A1(N7349), .S(n3881), .Z(n15467) );
  CMXI2X1 U26758 ( .A0(n15467), .A1(n15461), .S(n4142), .Z(n15474) );
  CMX2X1 U26759 ( .A0(n15462), .A1(n15474), .S(n3793), .Z(n15490) );
  CMXI2X1 U26760 ( .A0(n15463), .A1(n15490), .S(n3386), .Z(N9195) );
  CMX2X1 U26761 ( .A0(N7349), .A1(N7348), .S(n3862), .Z(n15470) );
  CMXI2X1 U26762 ( .A0(n15470), .A1(n15464), .S(n4142), .Z(n15480) );
  CMX2X1 U26763 ( .A0(n15465), .A1(n15480), .S(n3794), .Z(n15493) );
  CMXI2X1 U26764 ( .A0(n15466), .A1(n15493), .S(n3386), .Z(N9196) );
  CMX2X1 U26765 ( .A0(N7348), .A1(N7347), .S(n3869), .Z(n15473) );
  CMXI2X1 U26766 ( .A0(n15473), .A1(n15467), .S(n4142), .Z(n15483) );
  CMX2X1 U26767 ( .A0(n15468), .A1(n15483), .S(n3795), .Z(n15496) );
  CMXI2X1 U26768 ( .A0(n15469), .A1(n15496), .S(n3386), .Z(N9197) );
  CMX2X1 U26769 ( .A0(N7347), .A1(N7346), .S(n3870), .Z(n15479) );
  CMXI2X1 U26770 ( .A0(n15479), .A1(n15470), .S(n4142), .Z(n15486) );
  CMX2X1 U26771 ( .A0(n15471), .A1(n15486), .S(n3796), .Z(n15499) );
  CMXI2X1 U26772 ( .A0(n15472), .A1(n15499), .S(n3386), .Z(N9198) );
  CMX2X1 U26773 ( .A0(N7346), .A1(N7345), .S(n3871), .Z(n15482) );
  CMXI2X1 U26774 ( .A0(n15482), .A1(n15473), .S(n4142), .Z(n15489) );
  CMX2X1 U26775 ( .A0(n15474), .A1(n15489), .S(n3797), .Z(n15502) );
  CMXI2X1 U26776 ( .A0(n15475), .A1(n15502), .S(n3386), .Z(N9199) );
  CMX2X1 U26777 ( .A0(n15477), .A1(n15476), .S(n3805), .Z(n15728) );
  CMXI2X1 U26778 ( .A0(n15478), .A1(n15728), .S(n3386), .Z(N8371) );
  CMX2X1 U26779 ( .A0(N7345), .A1(N7344), .S(n3872), .Z(n15485) );
  CMXI2X1 U26780 ( .A0(n15485), .A1(n15479), .S(n4142), .Z(n15492) );
  CMX2X1 U26781 ( .A0(n15480), .A1(n15492), .S(n3806), .Z(n15505) );
  CMXI2X1 U26782 ( .A0(n15481), .A1(n15505), .S(n3386), .Z(N9200) );
  CMX2X1 U26783 ( .A0(N7344), .A1(N7343), .S(n3867), .Z(n15488) );
  CMXI2X1 U26784 ( .A0(n15488), .A1(n15482), .S(n4142), .Z(n15495) );
  CMX2X1 U26785 ( .A0(n15483), .A1(n15495), .S(n3775), .Z(n15508) );
  CMXI2X1 U26786 ( .A0(n15484), .A1(n15508), .S(n3386), .Z(N9201) );
  CMX2X1 U26787 ( .A0(N7343), .A1(N7342), .S(n3868), .Z(n15491) );
  CMXI2X1 U26788 ( .A0(n15491), .A1(n15485), .S(n4142), .Z(n15498) );
  CMX2X1 U26789 ( .A0(n15486), .A1(n15498), .S(n3810), .Z(n15513) );
  CMXI2X1 U26790 ( .A0(n15487), .A1(n15513), .S(n3386), .Z(N9202) );
  CMX2X1 U26791 ( .A0(N7342), .A1(N7341), .S(n3869), .Z(n15494) );
  CMXI2X1 U26792 ( .A0(n15494), .A1(n15488), .S(n4142), .Z(n15501) );
  CMX2X1 U26793 ( .A0(n15489), .A1(n15501), .S(n3796), .Z(n15516) );
  CMXI2X1 U26794 ( .A0(n15490), .A1(n15516), .S(n3386), .Z(N9203) );
  CMX2X1 U26795 ( .A0(N7341), .A1(N7340), .S(n3870), .Z(n15497) );
  CMXI2X1 U26796 ( .A0(n15497), .A1(n15491), .S(n4142), .Z(n15504) );
  CMX2X1 U26797 ( .A0(n15492), .A1(n15504), .S(n3797), .Z(n15519) );
  CMXI2X1 U26798 ( .A0(n15493), .A1(n15519), .S(n3385), .Z(N9204) );
  CMX2X1 U26799 ( .A0(N7340), .A1(N7339), .S(n3863), .Z(n15500) );
  CMXI2X1 U26800 ( .A0(n15500), .A1(n15494), .S(n4142), .Z(n15507) );
  CMX2X1 U26801 ( .A0(n15495), .A1(n15507), .S(n3805), .Z(n15522) );
  CMXI2X1 U26802 ( .A0(n15496), .A1(n15522), .S(n3389), .Z(N9205) );
  CMX2X1 U26803 ( .A0(N7339), .A1(N7338), .S(n3863), .Z(n15503) );
  CMXI2X1 U26804 ( .A0(n15503), .A1(n15497), .S(n4142), .Z(n15512) );
  CMX2X1 U26805 ( .A0(n15498), .A1(n15512), .S(n3806), .Z(n15525) );
  CMXI2X1 U26806 ( .A0(n15499), .A1(n15525), .S(n3389), .Z(N9206) );
  CMX2X1 U26807 ( .A0(N7338), .A1(N7337), .S(n3864), .Z(n15506) );
  CMXI2X1 U26808 ( .A0(n15506), .A1(n15500), .S(n4142), .Z(n15515) );
  CMX2X1 U26809 ( .A0(n15501), .A1(n15515), .S(n3807), .Z(n15528) );
  CMXI2X1 U26810 ( .A0(n15502), .A1(n15528), .S(n3389), .Z(N9207) );
  CMX2X1 U26811 ( .A0(N7337), .A1(N7336), .S(n3865), .Z(n15511) );
  CMXI2X1 U26812 ( .A0(n15511), .A1(n15503), .S(n4141), .Z(n15518) );
  CMX2X1 U26813 ( .A0(n15504), .A1(n15518), .S(n3794), .Z(n15531) );
  CMXI2X1 U26814 ( .A0(n15505), .A1(n15531), .S(n3388), .Z(N9208) );
  CMX2X1 U26815 ( .A0(N7336), .A1(N7335), .S(n3866), .Z(n15514) );
  CMXI2X1 U26816 ( .A0(n15514), .A1(n15506), .S(n4141), .Z(n15521) );
  CMX2X1 U26817 ( .A0(n15507), .A1(n15521), .S(n3807), .Z(n15534) );
  CMXI2X1 U26818 ( .A0(n15508), .A1(n15534), .S(n3388), .Z(N9209) );
  CMXI2X1 U26819 ( .A0(n15510), .A1(n15509), .S(n3388), .Z(N8372) );
  CMX2X1 U26820 ( .A0(N7335), .A1(N7334), .S(n3867), .Z(n15517) );
  CMXI2X1 U26821 ( .A0(n15517), .A1(n15511), .S(n4141), .Z(n15524) );
  CMX2X1 U26822 ( .A0(n15512), .A1(n15524), .S(n3808), .Z(n15537) );
  CMXI2X1 U26823 ( .A0(n15513), .A1(n15537), .S(n3388), .Z(N9210) );
  CMX2X1 U26824 ( .A0(N7334), .A1(N7333), .S(n3868), .Z(n15520) );
  CMXI2X1 U26825 ( .A0(n15520), .A1(n15514), .S(n4141), .Z(n15527) );
  CMX2X1 U26826 ( .A0(n15515), .A1(n15527), .S(n3809), .Z(n15540) );
  CMXI2X1 U26827 ( .A0(n15516), .A1(n15540), .S(n3388), .Z(N9211) );
  CMX2X1 U26828 ( .A0(N7333), .A1(N7332), .S(n3869), .Z(n15523) );
  CMXI2X1 U26829 ( .A0(n15523), .A1(n15517), .S(n4141), .Z(n15530) );
  CMX2X1 U26830 ( .A0(n15518), .A1(n15530), .S(n3810), .Z(n15545) );
  CMXI2X1 U26831 ( .A0(n15519), .A1(n15545), .S(n3388), .Z(N9212) );
  CMX2X1 U26832 ( .A0(N7332), .A1(N7331), .S(n3874), .Z(n15526) );
  CMXI2X1 U26833 ( .A0(n15526), .A1(n15520), .S(n4141), .Z(n15533) );
  CMX2X1 U26834 ( .A0(n15521), .A1(n15533), .S(n3811), .Z(n15548) );
  CMXI2X1 U26835 ( .A0(n15522), .A1(n15548), .S(n3388), .Z(N9213) );
  CMX2X1 U26836 ( .A0(N7331), .A1(N7330), .S(n3875), .Z(n15529) );
  CMXI2X1 U26837 ( .A0(n15529), .A1(n15523), .S(n4141), .Z(n15536) );
  CMX2X1 U26838 ( .A0(n15524), .A1(n15536), .S(n3812), .Z(n15551) );
  CMXI2X1 U26839 ( .A0(n15525), .A1(n15551), .S(n3388), .Z(N9214) );
  CMX2X1 U26840 ( .A0(N7330), .A1(N7329), .S(n3870), .Z(n15532) );
  CMXI2X1 U26841 ( .A0(n15532), .A1(n15526), .S(n4141), .Z(n15539) );
  CMX2X1 U26842 ( .A0(n15527), .A1(n15539), .S(n4306), .Z(n15554) );
  CMXI2X1 U26843 ( .A0(n15528), .A1(n15554), .S(n3388), .Z(N9215) );
  CMX2X1 U26844 ( .A0(N7329), .A1(N7328), .S(n3871), .Z(n15535) );
  CMXI2X1 U26845 ( .A0(n15535), .A1(n15529), .S(n4141), .Z(n15544) );
  CMX2X1 U26846 ( .A0(n15530), .A1(n15544), .S(n3771), .Z(n15557) );
  CMXI2X1 U26847 ( .A0(n15531), .A1(n15557), .S(n3388), .Z(N9216) );
  CMX2X1 U26848 ( .A0(N7328), .A1(N7327), .S(n3873), .Z(n15538) );
  CMXI2X1 U26849 ( .A0(n15538), .A1(n15532), .S(n4141), .Z(n15547) );
  CMX2X1 U26850 ( .A0(n15533), .A1(n15547), .S(n3772), .Z(n15560) );
  CMXI2X1 U26851 ( .A0(n15534), .A1(n15560), .S(n3388), .Z(N9217) );
  CMX2X1 U26852 ( .A0(N7327), .A1(N7326), .S(n3874), .Z(n15543) );
  CMXI2X1 U26853 ( .A0(n15543), .A1(n15535), .S(n4141), .Z(n15550) );
  CMX2X1 U26854 ( .A0(n15536), .A1(n15550), .S(n3773), .Z(n15563) );
  CMXI2X1 U26855 ( .A0(n15537), .A1(n15563), .S(n3387), .Z(N9218) );
  CMX2X1 U26856 ( .A0(N7326), .A1(N7325), .S(n3875), .Z(n15546) );
  CMXI2X1 U26857 ( .A0(n15546), .A1(n15538), .S(n4141), .Z(n15553) );
  CMX2X1 U26858 ( .A0(n15539), .A1(n15553), .S(n3774), .Z(n15566) );
  CMXI2X1 U26859 ( .A0(n15540), .A1(n15566), .S(n3387), .Z(N9219) );
  CMXI2X1 U26860 ( .A0(n15542), .A1(n15541), .S(n3387), .Z(N8373) );
  CMX2X1 U26861 ( .A0(N7325), .A1(N7324), .S(n3876), .Z(n15549) );
  CMXI2X1 U26862 ( .A0(n15549), .A1(n15543), .S(n4141), .Z(n15556) );
  CMX2X1 U26863 ( .A0(n15544), .A1(n15556), .S(n3775), .Z(n15569) );
  CMXI2X1 U26864 ( .A0(n15545), .A1(n15569), .S(n3387), .Z(N9220) );
  CMX2X1 U26865 ( .A0(N7324), .A1(N7323), .S(n3871), .Z(n15552) );
  CMXI2X1 U26866 ( .A0(n15552), .A1(n15546), .S(n4141), .Z(n15559) );
  CMX2X1 U26867 ( .A0(n15547), .A1(n15559), .S(n3776), .Z(n15572) );
  CMXI2X1 U26868 ( .A0(n15548), .A1(n15572), .S(n3390), .Z(N9221) );
  CMX2X1 U26869 ( .A0(N7323), .A1(N7322), .S(n3872), .Z(n15555) );
  CMXI2X1 U26870 ( .A0(n15555), .A1(n15549), .S(n4141), .Z(n15562) );
  CMX2X1 U26871 ( .A0(n15550), .A1(n15562), .S(n3777), .Z(n15577) );
  CMXI2X1 U26872 ( .A0(n15551), .A1(n15577), .S(n3390), .Z(N9222) );
  CMX2X1 U26873 ( .A0(N7322), .A1(N7321), .S(n3873), .Z(n15558) );
  CMXI2X1 U26874 ( .A0(n15558), .A1(n15552), .S(n4141), .Z(n15565) );
  CMX2X1 U26875 ( .A0(n15553), .A1(n15565), .S(n3794), .Z(n15580) );
  CMXI2X1 U26876 ( .A0(n15554), .A1(n15580), .S(n3390), .Z(N9223) );
  CMX2X1 U26877 ( .A0(N7321), .A1(N7320), .S(n3874), .Z(n15561) );
  CMXI2X1 U26878 ( .A0(n15561), .A1(n15555), .S(n4140), .Z(n15568) );
  CMX2X1 U26879 ( .A0(n15556), .A1(n15568), .S(n3792), .Z(n15583) );
  CMXI2X1 U26880 ( .A0(n15557), .A1(n15583), .S(n3390), .Z(N9224) );
  CMX2X1 U26881 ( .A0(N7320), .A1(N7319), .S(n3864), .Z(n15564) );
  CMXI2X1 U26882 ( .A0(n15564), .A1(n15558), .S(n4140), .Z(n15571) );
  CMX2X1 U26883 ( .A0(n15559), .A1(n15571), .S(n3793), .Z(n15586) );
  CMXI2X1 U26884 ( .A0(n15560), .A1(n15586), .S(n3390), .Z(N9225) );
  CMX2X1 U26885 ( .A0(N7319), .A1(N7318), .S(n3872), .Z(n15567) );
  CMXI2X1 U26886 ( .A0(n15567), .A1(n15561), .S(n4140), .Z(n15576) );
  CMX2X1 U26887 ( .A0(n15562), .A1(n15576), .S(n3794), .Z(n15589) );
  CMXI2X1 U26888 ( .A0(n15563), .A1(n15589), .S(n3390), .Z(N9226) );
  CMX2X1 U26889 ( .A0(N7318), .A1(N7317), .S(n3873), .Z(n15570) );
  CMXI2X1 U26890 ( .A0(n15570), .A1(n15564), .S(n4140), .Z(n15579) );
  CMX2X1 U26891 ( .A0(n15565), .A1(n15579), .S(n3795), .Z(n15592) );
  CMXI2X1 U26892 ( .A0(n15566), .A1(n15592), .S(n3390), .Z(N9227) );
  CMX2X1 U26893 ( .A0(N7317), .A1(N7316), .S(n3874), .Z(n15575) );
  CMXI2X1 U26894 ( .A0(n15575), .A1(n15567), .S(n4140), .Z(n15582) );
  CMX2X1 U26895 ( .A0(n15568), .A1(n15582), .S(n3796), .Z(n15595) );
  CMXI2X1 U26896 ( .A0(n15569), .A1(n15595), .S(n3390), .Z(N9228) );
  CMX2X1 U26897 ( .A0(N7316), .A1(N7315), .S(n3875), .Z(n15578) );
  CMXI2X1 U26898 ( .A0(n15578), .A1(n15570), .S(n4140), .Z(n15585) );
  CMX2X1 U26899 ( .A0(n15571), .A1(n15585), .S(n3797), .Z(n15598) );
  CMXI2X1 U26900 ( .A0(n15572), .A1(n15598), .S(n3390), .Z(N9229) );
  CMXI2X1 U26901 ( .A0(n15574), .A1(n15573), .S(n3390), .Z(N8374) );
  CMX2X1 U26902 ( .A0(N7315), .A1(N7314), .S(n3876), .Z(n15581) );
  CMXI2X1 U26903 ( .A0(n15581), .A1(n15575), .S(n4140), .Z(n15588) );
  CMX2X1 U26904 ( .A0(n15576), .A1(n15588), .S(n3805), .Z(n15601) );
  CMXI2X1 U26905 ( .A0(n15577), .A1(n15601), .S(n3389), .Z(N9230) );
  CMX2X1 U26906 ( .A0(N7314), .A1(N7313), .S(n3877), .Z(n15584) );
  CMXI2X1 U26907 ( .A0(n15584), .A1(n15578), .S(n4140), .Z(n15591) );
  CMX2X1 U26908 ( .A0(n15579), .A1(n15591), .S(n3806), .Z(n15604) );
  CMXI2X1 U26909 ( .A0(n15580), .A1(n15604), .S(n3389), .Z(N9231) );
  CMX2X1 U26910 ( .A0(N7313), .A1(N7312), .S(n3878), .Z(n15587) );
  CMXI2X1 U26911 ( .A0(n15587), .A1(n15581), .S(n4140), .Z(n15594) );
  CMX2X1 U26912 ( .A0(n15582), .A1(n15594), .S(n3807), .Z(n15609) );
  CMXI2X1 U26913 ( .A0(n15583), .A1(n15609), .S(n3389), .Z(N9232) );
  CMX2X1 U26914 ( .A0(N7312), .A1(N7311), .S(n3876), .Z(n15590) );
  CMXI2X1 U26915 ( .A0(n15590), .A1(n15584), .S(n4140), .Z(n15597) );
  CMX2X1 U26916 ( .A0(n15585), .A1(n15597), .S(n3808), .Z(n15612) );
  CMXI2X1 U26917 ( .A0(n15586), .A1(n15612), .S(n3389), .Z(N9233) );
  CMX2X1 U26918 ( .A0(N7311), .A1(N7310), .S(n3877), .Z(n15593) );
  CMXI2X1 U26919 ( .A0(n15593), .A1(n15587), .S(n4140), .Z(n15600) );
  CMX2X1 U26920 ( .A0(n15588), .A1(n15600), .S(n3809), .Z(n15615) );
  CMXI2X1 U26921 ( .A0(n15589), .A1(n15615), .S(n3389), .Z(N9234) );
  CMX2X1 U26922 ( .A0(N7310), .A1(N7309), .S(n3879), .Z(n15596) );
  CMXI2X1 U26923 ( .A0(n15596), .A1(n15590), .S(n4140), .Z(n15603) );
  CMX2X1 U26924 ( .A0(n15591), .A1(n15603), .S(n3810), .Z(n15618) );
  CMXI2X1 U26925 ( .A0(n15592), .A1(n15618), .S(n3389), .Z(N9235) );
  CMX2X1 U26926 ( .A0(N7309), .A1(N7308), .S(n3880), .Z(n15599) );
  CMXI2X1 U26927 ( .A0(n15599), .A1(n15593), .S(n4140), .Z(n15608) );
  CMX2X1 U26928 ( .A0(n15594), .A1(n15608), .S(n3811), .Z(n15621) );
  CMXI2X1 U26929 ( .A0(n15595), .A1(n15621), .S(n3389), .Z(N9236) );
  CMX2X1 U26930 ( .A0(N7308), .A1(N7307), .S(n3877), .Z(n15602) );
  CMXI2X1 U26931 ( .A0(n15602), .A1(n15596), .S(n4140), .Z(n15611) );
  CMX2X1 U26932 ( .A0(n15597), .A1(n15611), .S(n3812), .Z(n15624) );
  CMXI2X1 U26933 ( .A0(n15598), .A1(n15624), .S(n3389), .Z(N9237) );
  CMX2X1 U26934 ( .A0(N7307), .A1(N7306), .S(n3878), .Z(n15607) );
  CMXI2X1 U26935 ( .A0(n15607), .A1(n15599), .S(n4140), .Z(n15614) );
  CMX2X1 U26936 ( .A0(n15600), .A1(n15614), .S(n4306), .Z(n15627) );
  CMXI2X1 U26937 ( .A0(n15601), .A1(n15627), .S(n3392), .Z(N9238) );
  CMX2X1 U26938 ( .A0(N7306), .A1(N7305), .S(n3879), .Z(n15610) );
  CMXI2X1 U26939 ( .A0(n15610), .A1(n15602), .S(n4140), .Z(n15617) );
  CMX2X1 U26940 ( .A0(n15603), .A1(n15617), .S(n3771), .Z(n15630) );
  CMXI2X1 U26941 ( .A0(n15604), .A1(n15630), .S(n3392), .Z(N9239) );
  CMXI2X1 U26942 ( .A0(n15606), .A1(n15605), .S(n3392), .Z(N8375) );
  CMX2X1 U26943 ( .A0(N7305), .A1(N7304), .S(n3880), .Z(n15613) );
  CMXI2X1 U26944 ( .A0(n15613), .A1(n15607), .S(n4139), .Z(n15620) );
  CMX2X1 U26945 ( .A0(n15608), .A1(n15620), .S(n3791), .Z(n15633) );
  CMXI2X1 U26946 ( .A0(n15609), .A1(n15633), .S(n3392), .Z(N9240) );
  CMX2X1 U26947 ( .A0(N7304), .A1(N7303), .S(n3875), .Z(n15616) );
  CMXI2X1 U26948 ( .A0(n15616), .A1(n15610), .S(n4139), .Z(n15623) );
  CMX2X1 U26949 ( .A0(n15611), .A1(n15623), .S(n3792), .Z(n15636) );
  CMXI2X1 U26950 ( .A0(n15612), .A1(n15636), .S(n3392), .Z(N9241) );
  CMX2X1 U26951 ( .A0(N7303), .A1(N7302), .S(n3876), .Z(n15619) );
  CMXI2X1 U26952 ( .A0(n15619), .A1(n15613), .S(n4139), .Z(n15626) );
  CMX2X1 U26953 ( .A0(n15614), .A1(n15626), .S(n3793), .Z(n15641) );
  CMXI2X1 U26954 ( .A0(n15615), .A1(n15641), .S(n3392), .Z(N9242) );
  CMX2X1 U26955 ( .A0(N7302), .A1(N7301), .S(n3877), .Z(n15622) );
  CMXI2X1 U26956 ( .A0(n15622), .A1(n15616), .S(n4139), .Z(n15629) );
  CMX2X1 U26957 ( .A0(n15617), .A1(n15629), .S(n3794), .Z(n15644) );
  CMXI2X1 U26958 ( .A0(n15618), .A1(n15644), .S(n3391), .Z(N9243) );
  CMX2X1 U26959 ( .A0(N7301), .A1(N7300), .S(n3878), .Z(n15625) );
  CMXI2X1 U26960 ( .A0(n15625), .A1(n15619), .S(n4139), .Z(n15632) );
  CMX2X1 U26961 ( .A0(n15620), .A1(n15632), .S(n3795), .Z(n15647) );
  CMXI2X1 U26962 ( .A0(n15621), .A1(n15647), .S(n3391), .Z(N9244) );
  CMX2X1 U26963 ( .A0(N7300), .A1(N7299), .S(n3865), .Z(n15628) );
  CMXI2X1 U26964 ( .A0(n15628), .A1(n15622), .S(n4139), .Z(n15635) );
  CMX2X1 U26965 ( .A0(n15623), .A1(n15635), .S(n3796), .Z(n15650) );
  CMXI2X1 U26966 ( .A0(n15624), .A1(n15650), .S(n3391), .Z(N9245) );
  CMX2X1 U26967 ( .A0(N7299), .A1(N7298), .S(n3881), .Z(n15631) );
  CMXI2X1 U26968 ( .A0(n15631), .A1(n15625), .S(n4139), .Z(n15640) );
  CMX2X1 U26969 ( .A0(n15626), .A1(n15640), .S(n3797), .Z(n15653) );
  CMXI2X1 U26970 ( .A0(n15627), .A1(n15653), .S(n3391), .Z(N9246) );
  CMX2X1 U26971 ( .A0(N7298), .A1(N7297), .S(n3862), .Z(n15634) );
  CMXI2X1 U26972 ( .A0(n15634), .A1(n15628), .S(n4139), .Z(n15643) );
  CMX2X1 U26973 ( .A0(n15629), .A1(n15643), .S(n3805), .Z(n15656) );
  CMXI2X1 U26974 ( .A0(n15630), .A1(n15656), .S(n3391), .Z(N9247) );
  CMX2X1 U26975 ( .A0(N7297), .A1(N7296), .S(n3863), .Z(n15639) );
  CMXI2X1 U26976 ( .A0(n15639), .A1(n15631), .S(n4139), .Z(n15646) );
  CMX2X1 U26977 ( .A0(n15632), .A1(n15646), .S(n3806), .Z(n15659) );
  CMXI2X1 U26978 ( .A0(n15633), .A1(n15659), .S(n3391), .Z(N9248) );
  CMX2X1 U26979 ( .A0(N7296), .A1(N7295), .S(n3864), .Z(n15642) );
  CMXI2X1 U26980 ( .A0(n15642), .A1(n15634), .S(n4139), .Z(n15649) );
  CMX2X1 U26981 ( .A0(n15635), .A1(n15649), .S(n3809), .Z(n15662) );
  CMXI2X1 U26982 ( .A0(n15636), .A1(n15662), .S(n3391), .Z(N9249) );
  CMXI2X1 U26983 ( .A0(n15638), .A1(n15637), .S(n3391), .Z(N8376) );
  CMX2X1 U26984 ( .A0(N7295), .A1(N7294), .S(n3865), .Z(n15645) );
  CMXI2X1 U26985 ( .A0(n15645), .A1(n15639), .S(n4139), .Z(n15652) );
  CMX2X1 U26986 ( .A0(n15640), .A1(n15652), .S(n3794), .Z(n15665) );
  CMXI2X1 U26987 ( .A0(n15641), .A1(n15665), .S(n3391), .Z(N9250) );
  CMX2X1 U26988 ( .A0(N7294), .A1(N7293), .S(n3866), .Z(n15648) );
  CMXI2X1 U26989 ( .A0(n15648), .A1(n15642), .S(n4139), .Z(n15655) );
  CMX2X1 U26990 ( .A0(n15643), .A1(n15655), .S(n3806), .Z(n15668) );
  CMXI2X1 U26991 ( .A0(n15644), .A1(n15668), .S(n3391), .Z(N9251) );
  CMX2X1 U26992 ( .A0(N7293), .A1(N7292), .S(n3867), .Z(n15651) );
  CMXI2X1 U26993 ( .A0(n15651), .A1(n15645), .S(n4139), .Z(n15658) );
  CMX2X1 U26994 ( .A0(n15646), .A1(n15658), .S(n3807), .Z(n15673) );
  CMXI2X1 U26995 ( .A0(n15647), .A1(n15673), .S(n3391), .Z(N9252) );
  CMX2X1 U26996 ( .A0(N7292), .A1(N7291), .S(n3878), .Z(n15654) );
  CMXI2X1 U26997 ( .A0(n15654), .A1(n15648), .S(n4139), .Z(n15661) );
  CMX2X1 U26998 ( .A0(n15649), .A1(n15661), .S(n3808), .Z(n15676) );
  CMXI2X1 U26999 ( .A0(n15650), .A1(n15676), .S(n3390), .Z(N9253) );
  CMX2X1 U27000 ( .A0(N7291), .A1(N7290), .S(n3879), .Z(n15657) );
  CMXI2X1 U27001 ( .A0(n15657), .A1(n15651), .S(n4139), .Z(n15664) );
  CMX2X1 U27002 ( .A0(n15652), .A1(n15664), .S(n3809), .Z(n15679) );
  CMXI2X1 U27003 ( .A0(n15653), .A1(n15679), .S(n3394), .Z(N9254) );
  CMX2X1 U27004 ( .A0(N7290), .A1(N7289), .S(n3868), .Z(n15660) );
  CMXI2X1 U27005 ( .A0(n15660), .A1(n15654), .S(n4139), .Z(n15667) );
  CMX2X1 U27006 ( .A0(n15655), .A1(n15667), .S(n3810), .Z(n15682) );
  CMXI2X1 U27007 ( .A0(n15656), .A1(n15682), .S(n3394), .Z(N9255) );
  CMX2X1 U27008 ( .A0(N7289), .A1(N7288), .S(n3869), .Z(n15663) );
  CMXI2X1 U27009 ( .A0(n15663), .A1(n15657), .S(n4138), .Z(n15672) );
  CMX2X1 U27010 ( .A0(n15658), .A1(n15672), .S(n3773), .Z(n15685) );
  CMXI2X1 U27011 ( .A0(n15659), .A1(n15685), .S(n3393), .Z(N9256) );
  CMX2X1 U27012 ( .A0(N7288), .A1(N7287), .S(n3881), .Z(n15666) );
  CMXI2X1 U27013 ( .A0(n15666), .A1(n15660), .S(n4138), .Z(n15675) );
  CMX2X1 U27014 ( .A0(n15661), .A1(n15675), .S(n3807), .Z(n15688) );
  CMXI2X1 U27015 ( .A0(n15662), .A1(n15688), .S(n3393), .Z(N9257) );
  CMX2X1 U27016 ( .A0(N7287), .A1(N7286), .S(n3862), .Z(n15671) );
  CMXI2X1 U27017 ( .A0(n15671), .A1(n15663), .S(n4138), .Z(n15678) );
  CMX2X1 U27018 ( .A0(n15664), .A1(n15678), .S(n3808), .Z(n15692) );
  CMXI2X1 U27019 ( .A0(n15665), .A1(n15692), .S(n3393), .Z(N9258) );
  CMX2X1 U27020 ( .A0(N7286), .A1(N7285), .S(n3863), .Z(n15674) );
  CMXI2X1 U27021 ( .A0(n15674), .A1(n15666), .S(n4138), .Z(n15681) );
  CMX2X1 U27022 ( .A0(n15667), .A1(n15681), .S(n3809), .Z(n15696) );
  CMXI2X1 U27023 ( .A0(n15668), .A1(n15696), .S(n3393), .Z(N9259) );
  CMXI2X1 U27024 ( .A0(n15670), .A1(n15669), .S(n3393), .Z(N8377) );
  CMXI2X1 U27025 ( .A0(n15677), .A1(n15671), .S(n4138), .Z(n15684) );
  CMX2X1 U27026 ( .A0(n15672), .A1(n15684), .S(n3810), .Z(n15699) );
  CMXI2X1 U27027 ( .A0(n15673), .A1(n15699), .S(n3393), .Z(N9260) );
  CMX2X1 U27028 ( .A0(N7284), .A1(N7283), .S(n3879), .Z(n15680) );
  CMXI2X1 U27029 ( .A0(n15680), .A1(n15674), .S(n4138), .Z(n15687) );
  CMX2X1 U27030 ( .A0(n15675), .A1(n15687), .S(n3811), .Z(n15702) );
  CMXI2X1 U27031 ( .A0(n15676), .A1(n15702), .S(n3393), .Z(N9261) );
  CMX2X1 U27032 ( .A0(N7283), .A1(N7282), .S(n3880), .Z(n15683) );
  CMXI2X1 U27033 ( .A0(n15683), .A1(n15677), .S(n4138), .Z(n15691) );
  CMX2X1 U27034 ( .A0(n15678), .A1(n15691), .S(n3812), .Z(n15707) );
  CMXI2X1 U27035 ( .A0(n15679), .A1(n15707), .S(n3393), .Z(N9262) );
  CMX2X1 U27036 ( .A0(N7282), .A1(N7281), .S(n3878), .Z(n15686) );
  CMXI2X1 U27037 ( .A0(n15686), .A1(n15680), .S(n4138), .Z(n15695) );
  CMX2X1 U27038 ( .A0(n15681), .A1(n15695), .S(n4306), .Z(n15710) );
  CMXI2X1 U27039 ( .A0(n15682), .A1(n15710), .S(n3393), .Z(N9263) );
  CMXI2X1 U27040 ( .A0(n15689), .A1(n15683), .S(n4138), .Z(n15698) );
  CMX2X1 U27041 ( .A0(n15684), .A1(n15698), .S(n3771), .Z(n15712) );
  CMXI2X1 U27042 ( .A0(n15685), .A1(n15712), .S(n3393), .Z(N9264) );
  CMXI2X1 U27043 ( .A0(n15693), .A1(n15686), .S(n4138), .Z(n15701) );
  CMX2X1 U27044 ( .A0(n15687), .A1(n15701), .S(n3772), .Z(n15714) );
  CMXI2X1 U27045 ( .A0(n15688), .A1(n15714), .S(n3393), .Z(N9265) );
  CMXI2X1 U27046 ( .A0(n15690), .A1(n15689), .S(n4138), .Z(n15706) );
  CMX2X1 U27047 ( .A0(n15691), .A1(n15706), .S(n3773), .Z(n15716) );
  CMXI2X1 U27048 ( .A0(n15692), .A1(n15716), .S(n3392), .Z(N9266) );
  CMXI2X1 U27049 ( .A0(n15694), .A1(n15693), .S(n4138), .Z(n15709) );
  CMX2X1 U27050 ( .A0(n15695), .A1(n15709), .S(n3774), .Z(n15718) );
  CMXI2X1 U27051 ( .A0(n15696), .A1(n15718), .S(n3392), .Z(N9267) );
  CMX2X1 U27052 ( .A0(n15698), .A1(n15697), .S(n3775), .Z(n15720) );
  CMXI2X1 U27053 ( .A0(n15699), .A1(n15720), .S(n3392), .Z(N9268) );
  CMX2X1 U27054 ( .A0(n15701), .A1(n15700), .S(n3812), .Z(n15722) );
  CMXI2X1 U27055 ( .A0(n15702), .A1(n15722), .S(n3392), .Z(N9269) );
  CMXI2X1 U27056 ( .A0(n15704), .A1(n15703), .S(n3392), .Z(N8378) );
  CMX2X1 U27057 ( .A0(n15706), .A1(n15705), .S(n3771), .Z(n15724) );
  CMXI2X1 U27058 ( .A0(n15707), .A1(n15724), .S(n3355), .Z(N9270) );
  CMX2X1 U27059 ( .A0(n15709), .A1(n15708), .S(n3809), .Z(n15726) );
  CMXI2X1 U27060 ( .A0(n15710), .A1(n15726), .S(n3354), .Z(N9271) );
  CMXI2X1 U27061 ( .A0(n15712), .A1(n15711), .S(n3353), .Z(N9272) );
  CMXI2X1 U27062 ( .A0(n15714), .A1(n15713), .S(n3352), .Z(N9273) );
  CMXI2X1 U27063 ( .A0(n15716), .A1(n15715), .S(n3390), .Z(N9274) );
  CMXI2X1 U27064 ( .A0(n15718), .A1(n15717), .S(n3389), .Z(N9275) );
  CMXI2X1 U27065 ( .A0(n15720), .A1(n15719), .S(n3382), .Z(N9276) );
  CMXI2X1 U27066 ( .A0(n15722), .A1(n15721), .S(n3371), .Z(N9277) );
  CMXI2X1 U27067 ( .A0(n15724), .A1(n15723), .S(n3359), .Z(N9278) );
  CMXI2X1 U27068 ( .A0(n15726), .A1(n15725), .S(n3358), .Z(N9279) );
  CMXI2X1 U27069 ( .A0(n15728), .A1(n15727), .S(n3393), .Z(N8379) );
  CMXI2X1 U27070 ( .A0(n15730), .A1(n15729), .S(n3392), .Z(N8289) );
endmodule

